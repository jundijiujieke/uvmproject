module imdct_rom257x64(
clk,
en,
addr,

dout
);

input clk;
input en;
input [8:0] addr;

output reg [63:0] dout;

reg [63:0] mem[0:256]={ 
64'h40000000_00000000, 
64'h40323034_003243f1, 
64'h406438cf_006487c4, 
64'h409619b2_0096cb58, 
64'h40c7d2bd_00c90e90, 
64'h40f963d3_00fb514b, 
64'h412accd4_012d936c, 
64'h415c0da3_015fd4d2, 
64'h418d2621_0192155f, 
64'h41be162f_01c454f5, 
64'h41eeddaf_01f69373, 
64'h421f7c84_0228d0bb, 
64'h424ff28f_025b0caf, 
64'h42803fb2_028d472e, 
64'h42b063d0_02bf801a, 
64'h42e05ecb_02f1b755, 
64'h43103085_0323ecbe, 
64'h433fd8e1_03562038, 
64'h436f57c1_038851a2, 
64'h439ead09_03ba80df, 
64'h43cdd89a_03ecadcf, 
64'h43fcda59_041ed854, 
64'h442bb227_0451004d, 
64'h445a5fe8_0483259d, 
64'h4488e37f_04b54825, 
64'h44b73ccf_04e767c5, 
64'h44e56bbd_0519845e, 
64'h4513702a_054b9dd3, 
64'h454149fc_057db403, 
64'h456ef916_05afc6d0,
64'h459c7d5a_05e1d61b, 
64'h45c9d6af_0613e1c5, 
64'h45f704f7_0645e9af, 
64'h46240816_0677edbb, 
64'h4650dff1_06a9edc9, 
64'h467d8c6d_06dbe9bb, 
64'h46aa0d6d_070de172, 
64'h46d662d6_073fd4cf, 
64'h47028c8d_0771c3b3, 
64'h472e8a76_07a3adff, 
64'h475a5c77_07d59396, 
64'h47860275_08077457, 
64'h47b17c54_08395024, 
64'h47dcc9f9_086b26de, 
64'h4807eb4b_089cf867,
64'h4832e02d_08cec4a0, 
64'h485da887_09008b6a, 
64'h4888443d_09324ca7, 
64'h48b2b335_09640837, 
64'h48dcf556_0995bdfd, 
64'h49070a84_09c76dd8, 
64'h4930f2a6_09f917ac, 
64'h495aada2_0a2abb59, 
64'h49843b5f_0a5c58c0, 
64'h49ad9bc2_0a8defc3, 
64'h49d6ceb3_0abf8043, 
64'h49ffd417_0af10a22, 
64'h4a28abd6_0b228d42, 
64'h4a5155d6_0b540982, 
64'h4a79d1ff_0b857ec7, 
64'h4aa22036_0bb6ecef, 
64'h4aca4065_0be853de, 
64'h4af23270_0c19b374, 
64'h4b19f641_0c4b0b94, 
64'h4b418bbe_0c7c5c1e, 
64'h4b68f2cf_0cada4f5, 
64'h4b902b5c_0cdee5f9, 
64'h4bb7354d_0d101f0e, 
64'h4bde1089_0d415013, 
64'h4c04bcf8_0d7278eb, 
64'h4c2b3a84_0da39978, 
64'h4c518913_0dd4b19a, 
64'h4c77a88e_0e05c135, 
64'h4c9d98de_0e36c82a, 
64'h4cc359ec_0e67c65a, 
64'h4ce8eb9f_0e98bba7, 
64'h4d0e4de2_0ec9a7f3, 
64'h4d33809c_0efa8b20, 
64'h4d5883b7_0f2b650f, 
64'h4d7d571c_0f5c35a3, 
64'h4da1fab5_0f8cfcbe, 
64'h4dc66e6a_0fbdba40, 
64'h4deab226_0fee6e0d, 
64'h4e0ec5d1_101f1807, 
64'h4e32a956_104fb80e, 
64'h4e565c9f_10804e06, 
64'h4e79df95_10b0d9d0, 
64'h4e9d3222_10e15b4e, 
64'h4ec05432_1111d263, 
64'h4ee345ad_11423ef0, 
64'h4f06067f_1172a0d7, 
64'h4f289692_11a2f7fc, 
64'h4f4af5d1_11d3443f, 
64'h4f6d2427_12038584, 
64'h4f8f217e_1233bbac, 
64'h4fb0edc1_1263e699, 
64'h4fd288dc_1294062f, 
64'h4ff3f2bb_12c41a4f, 
64'h50152b47_12f422db, 
64'h5036326e_13241fb6, 
64'h50570819_135410c3, 
64'h5077ac37_1383f5e3, 
64'h50981eb1_13b3cefa, 
64'h50b85f74_13e39be9, 
64'h50d86e6d_14135c94, 
64'h50f84b87_144310dd, 
64'h5117f6ae_1472b8a5, 
64'h51376fd0_14a253d1, 
64'h5156b6d9_14d1e242, 
64'h5175cbb5_150163dc, 
64'h5194ae52_1530d881, 
64'h51b35e9b_15604013, 
64'h51d1dc80_158f9a76, 
64'h51f027eb_15bee78c, 
64'h520e40cc_15ee2738, 
64'h522c270f_161d595d, 
64'h5249daa2_164c7ddd, 
64'h52675b72_167b949d, 
64'h5284a96e_16aa9d7e, 
64'h52a1c482_16d99864, 
64'h52beac9f_17088531, 
64'h52db61b0_173763c9, 
64'h52f7e3a6_1766340f, 
64'h5314326d_1794f5e6, 
64'h53304df6_17c3a931, 
64'h534c362d_17f24dd3, 
64'h5367eb03_1820e3b0, 
64'h53836c66_184f6aab, 
64'h539eba45_187de2a7, 
64'h53b9d48f_18ac4b87, 
64'h53d4bb34_18daa52f, 
64'h53ef6e23_1908ef82, 
64'h5409ed4b_19372a64, 
64'h5424389d_196555b8, 
64'h543e5007_19937161, 
64'h5458337a_19c17d44, 
64'h5471e2e6_19ef7944, 
64'h548b5e3b_1a1d6544, 
64'h54a4a56a_1a4b4128, 
64'h54bdb862_1a790cd4, 
64'h54d69714_1aa6c82b, 
64'h54ef4171_1ad47312, 
64'h5507b76a_1b020d6c, 
64'h551ff8ef_1b2f971e, 
64'h553805f2_1b5d100a, 
64'h554fde64_1b8a7815, 
64'h55678236_1bb7cf23, 
64'h557ef15a_1be51518, 
64'h55962bc0_1c1249d8, 
64'h55ad315b_1c3f6d47, 
64'h55c4021d_1c6c7f4a, 
64'h55da9df7_1c997fc4, 
64'h55f104dc_1cc66e99, 
64'h560736bd_1cf34baf, 
64'h561d338d_1d2016e9, 
64'h5632fb3f_1d4cd02c, 
64'h56488dc5_1d79775c, 
64'h565deb11_1da60c5d, 
64'h56731317_1dd28f15, 
64'h568805c9_1dfeff67, 
64'h569cc31b_1e2b5d38, 
64'h56b14b00_1e57a86d, 
64'h56c59d6a_1e83e0eb, 
64'h56d9ba4e_1eb00696, 
64'h56eda1a0_1edc1953, 
64'h57015352_1f081907, 
64'h5714cf59_1f340596, 
64'h572815a8_1f5fdee6, 
64'h573b2635_1f8ba4dc, 
64'h574e00f2_1fb7575c, 
64'h5760a5d5_1fe2f64c, 
64'h577314d2_200e8190, 
64'h57854ddd_2039f90f, 
64'h579750ec_20655cac, 
64'h57a91df2_2090ac4d, 
64'h57bab4e6_20bbe7d8, 
64'h57cc15bc_20e70f32, 
64'h57dd406a_21122240, 
64'h57ee34e5_213d20e8, 
64'h57fef323_21680b0f, 
64'h580f7b19_2192e09b, 
64'h581fccbc_21bda171, 
64'h582fe804_21e84d76, 
64'h583fcce6_2212e492, 
64'h584f7b58_223d66a8, 
64'h585ef351_2267d3a0, 
64'h586e34c7_22922b5e, 
64'h587d3fb0_22bc6dca, 
64'h588c1404_22e69ac8, 
64'h589ab1b9_2310b23e, 
64'h58a918c6_233ab414, 
64'h58b74923_2364a02e, 
64'h58c542c5_238e7673, 
64'h58d305a6_23b836ca, 
64'h58e091bd_23e1e117, 
64'h58ede700_240b7543, 
64'h58fb0568_2434f332, 
64'h5907eced_245e5acc, 
64'h59149d87_2487abf7, 
64'h5921172e_24b0e699, 
64'h592d59da_24da0a9a, 
64'h59396584_250317df, 
64'h59453a24_252c0e4f, 
64'h5950d7b3_2554edd1, 
64'h595c3e2a_257db64c, 
64'h59676d82_25a667a7, 
64'h597265b4_25cf01c8, 
64'h597d26b8_25f78497, 
64'h5987b08a_261feffa, 
64'h59920321_264843d9, 
64'h599c1e78_2670801a, 
64'h59a60288_2698a4a6, 
64'h59afaf4c_26c0b162, 
64'h59b924bc_26e8a637, 
64'h59c262d5_2710830c, 
64'h59cb698f_273847c8, 
64'h59d438e5_275ff452, 
64'h59dcd0d3_27878893, 
64'h59e53151_27af0472, 
64'h59ed5a5c_27d667d5, 
64'h59f54bee_27fdb2a7, 
64'h59fd0603_2824e4cc, 
64'h5a048895_284bfe2f, 
64'h5a0bd3a1_2872feb6, 
64'h5a12e720_2899e64a, 
64'h5a19c310_28c0b4d2, 
64'h5a20676c_28e76a37, 
64'h5a26d42f_290e0661, 
64'h5a2d0957_29348937, 
64'h5a3306de_295af2a3, 
64'h5a38ccc2_2981428c, 
64'h5a3e5afe_29a778db, 
64'h5a43b190_29cd9578, 
64'h5a48d074_29f3984c, 
64'h5a4db7a6_2a19813f, 
64'h5a526725_2a3f503a, 
64'h5a56deec_2a650525, 
64'h5a5b1efa_2a8a9fea, 
64'h5a5f274b_2ab02071, 
64'h5a62f7dd_2ad586a3, 
64'h5a6690ae_2afad269, 
64'h5a69f1bb_2b2003ac, 
64'h5a6d1b03_2b451a55, 
64'h5a700c84_2b6a164d, 
64'h5a72c63b_2b8ef77d, 
64'h5a754827_2bb3bdce, 
64'h5a779246_2bd8692b, 
64'h5a79a498_2bfcf97c, 
64'h5a7b7f1a_2c216eaa, 
64'h5a7d21cc_2c45c8a0, 
64'h5a7e8cac_2c6a0746, 
64'h5a7fbfbb_2c8e2a87, 
64'h5a80baf6_2cb2324c, 
64'h5a817e5d_2cd61e7f, 
64'h5a8209f1_2cf9ef09, 
64'h5a825db0_2d1da3d5, 
64'h5a82799a_2d413ccd
};


always @(posedge clk) 
  if (en)
    dout <= mem[addr];

endmodule
