module rom_twidTabEven(
clk,
en,
addr,

dout
);

input clk;
input en;
input [9:0] addr;

output reg [31:0] dout;

reg [31:0] mem[0:503]={ 

32'h40000000,
32'h00000000,
32'h40000000,
32'h00000000,
32'h40000000,
32'h00000000,
32'h5a82799a,
32'hd2bec333,
32'h539eba45,
32'he7821d59,
32'h539eba45,
32'hc4df2862,
32'h40000000,
32'hc0000000,
32'h5a82799a,
32'hd2bec333,
32'h00000000,
32'hd2bec333,
32'h00000000,
32'hd2bec333,
32'h539eba45,
32'hc4df2862,
32'hac6145bb,
32'h187de2a7,
32'h40000000,
32'h00000000,
32'h40000000,
32'h00000000,
32'h40000000,
32'h00000000,
32'h4b418bbe,
32'hf383a3e2,
32'h45f704f7,
32'hf9ba1651,
32'h4fd288dc,
32'hed6bf9d1,
32'h539eba45,
32'he7821d59,
32'h4b418bbe,
32'hf383a3e2,
32'h58c542c5,
32'hdc71898d,
32'h58c542c5,
32'hdc71898d,
32'h4fd288dc,
32'hed6bf9d1,
32'h5a12e720,
32'hce86ff2a,
32'h5a82799a,
32'hd2bec333,
32'h539eba45,
32'he7821d59,
32'h539eba45,
32'hc4df2862,
32'h58c542c5,
32'hcac933ae,
32'h569cc31b,
32'he1d4a2c8,
32'h45f704f7,
32'hc04ee4b8,
32'h539eba45,
32'hc4df2862,
32'h58c542c5,
32'hdc71898d,
32'h3248d382,
32'hc13ad060,
32'h4b418bbe,
32'hc13ad060,
32'h5a12e720,
32'hd76619b6,
32'h1a4608ab,
32'hc78e9a1d,
32'h40000000,
32'hc0000000,
32'h5a82799a,
32'hd2bec333,
32'h00000000,
32'hd2bec333,
32'h3248d382,
32'hc13ad060,
32'h5a12e720,
32'hce86ff2a,
32'he5b9f755,
32'he1d4a2c8,
32'h22a2f4f8,
32'hc4df2862,
32'h58c542c5,
32'hcac933ae,
32'hcdb72c7e,
32'hf383a3e2,
32'h11a855df,
32'hcac933ae,
32'h569cc31b,
32'hc78e9a1d,
32'hba08fb09,
32'h0645e9af,
32'h00000000,
32'hd2bec333,
32'h539eba45,
32'hc4df2862,
32'hac6145bb,
32'h187de2a7,
32'hee57aa21,
32'hdc71898d,
32'h4fd288dc,
32'hc2c17d52,
32'ha5ed18e0,
32'h2899e64a,
32'hdd5d0b08,
32'he7821d59,
32'h4b418bbe,
32'hc13ad060,
32'ha73abd3b,
32'h3536cc52,
32'hcdb72c7e,
32'hf383a3e2,
32'h45f704f7,
32'hc04ee4b8,
32'hb02d7724,
32'h3d3e82ae,
32'h40000000,
32'h00000000,
32'h40000000,
32'h00000000,
32'h40000000,
32'h00000000,
32'h43103085,
32'hfcdc1342,
32'h418d2621,
32'hfe6deaa1,
32'h4488e37f,
32'hfb4ab7db,
32'h45f704f7,
32'hf9ba1651,
32'h43103085,
32'hfcdc1342,
32'h48b2b335,
32'hf69bf7c9,
32'h48b2b335,
32'hf69bf7c9,
32'h4488e37f,
32'hfb4ab7db,
32'h4c77a88e,
32'hf1fa3ecb,
32'h4b418bbe,
32'hf383a3e2,
32'h45f704f7,
32'hf9ba1651,
32'h4fd288dc,
32'hed6bf9d1,
32'h4da1fab5,
32'hf0730342,
32'h475a5c77,
32'hf82a6c6a,
32'h52beac9f,
32'he8f77acf,
32'h4fd288dc,
32'hed6bf9d1,
32'h48b2b335,
32'hf69bf7c9,
32'h553805f2,
32'he4a2eff6,
32'h51d1dc80,
32'hea70658a,
32'h49ffd417,
32'hf50ef5de,
32'h573b2635,
32'he0745b24,
32'h539eba45,
32'he7821d59,
32'h4b418bbe,
32'hf383a3e2,
32'h58c542c5,
32'hdc71898d,
32'h553805f2,
32'he4a2eff6,
32'h4c77a88e,
32'hf1fa3ecb,
32'h59d438e5,
32'hd8a00bae,
32'h569cc31b,
32'he1d4a2c8,
32'h4da1fab5,
32'hf0730342,
32'h5a6690ae,
32'hd5052d97,
32'h57cc15bc,
32'hdf18f0ce,
32'h4ec05432,
32'heeee2d9d,
32'h5a7b7f1a,
32'hd1a5ef90,
32'h58c542c5,
32'hdc71898d,
32'h4fd288dc,
32'hed6bf9d1,
32'h5a12e720,
32'hce86ff2a,
32'h5987b08a,
32'hd9e01006,
32'h50d86e6d,
32'hebeca36c,
32'h592d59da,
32'hcbacb0bf,
32'h5a12e720,
32'hd76619b6,
32'h51d1dc80,
32'hea70658a,
32'h57cc15bc,
32'hc91af976,
32'h5a6690ae,
32'hd5052d97,
32'h52beac9f,
32'he8f77acf,
32'h55f104dc,
32'hc6d569be,
32'h5a82799a,
32'hd2bec333,
32'h539eba45,
32'he7821d59,
32'h539eba45,
32'hc4df2862,
32'h5a6690ae,
32'hd09441bb,
32'h5471e2e6,
32'he61086bc,
32'h50d86e6d,
32'hc33aee27,
32'h5a12e720,
32'hce86ff2a,
32'h553805f2,
32'he4a2eff6,
32'h4da1fab5,
32'hc1eb0209,
32'h5987b08a,
32'hcc983f70,
32'h55f104dc,
32'he3399167,
32'h49ffd417,
32'hc0f1360b,
32'h58c542c5,
32'hcac933ae,
32'h569cc31b,
32'he1d4a2c8,
32'h45f704f7,
32'hc04ee4b8,
32'h57cc15bc,
32'hc91af976,
32'h573b2635,
32'he0745b24,
32'h418d2621,
32'hc004ef3f,
32'h569cc31b,
32'hc78e9a1d,
32'h57cc15bc,
32'hdf18f0ce,
32'h3cc85709,
32'hc013bc39,
32'h553805f2,
32'hc6250a18,
32'h584f7b58,
32'hddc29958,
32'h37af354c,
32'hc07b371e,
32'h539eba45,
32'hc4df2862,
32'h58c542c5,
32'hdc71898d,
32'h3248d382,
32'hc13ad060,
32'h51d1dc80,
32'hc3bdbdf6,
32'h592d59da,
32'hdb25f566,
32'h2c9caf6c,
32'hc2517e31,
32'h4fd288dc,
32'hc2c17d52,
32'h5987b08a,
32'hd9e01006,
32'h26b2a794,
32'hc3bdbdf6,
32'h4da1fab5,
32'hc1eb0209,
32'h59d438e5,
32'hd8a00bae,
32'h2092f05f,
32'hc57d965d,
32'h4b418bbe,
32'hc13ad060,
32'h5a12e720,
32'hd76619b6,
32'h1a4608ab,
32'hc78e9a1d,
32'h48b2b335,
32'hc0b15502,
32'h5a43b190,
32'hd6326a88,
32'h13d4ae08,
32'hc9edeb50,
32'h45f704f7,
32'hc04ee4b8,
32'h5a6690ae,
32'hd5052d97,
32'h0d47d096,
32'hcc983f70,
32'h43103085,
32'hc013bc39,
32'h5a7b7f1a,
32'hd3de9156,
32'h06a886a0,
32'hcf89e3e8,
32'h40000000,
32'hc0000000,
32'h5a82799a,
32'hd2bec333,
32'h00000000,
32'hd2bec333,
32'h3cc85709,
32'hc013bc39,
32'h5a7b7f1a,
32'hd1a5ef90,
32'hf9577960,
32'hd6326a88,
32'h396b3199,
32'hc04ee4b8,
32'h5a6690ae,
32'hd09441bb,
32'hf2b82f6a,
32'hd9e01006,
32'h35eaa2c7,
32'hc0b15502,
32'h5a43b190,
32'hcf89e3e8,
32'hec2b51f8,
32'hddc29958,
32'h3248d382,
32'hc13ad060,
32'h5a12e720,
32'hce86ff2a,
32'he5b9f755,
32'he1d4a2c8,
32'h2e88013a,
32'hc1eb0209,
32'h59d438e5,
32'hcd8bbb6d,
32'hdf6d0fa1,
32'he61086bc,
32'h2aaa7c7f,
32'hc2c17d52,
32'h5987b08a,
32'hcc983f70,
32'hd94d586c,
32'hea70658a,
32'h26b2a794,
32'hc3bdbdf6,
32'h592d59da,
32'hcbacb0bf,
32'hd3635094,
32'heeee2d9d,
32'h22a2f4f8,
32'hc4df2862,
32'h58c542c5,
32'hcac933ae,
32'hcdb72c7e,
32'hf383a3e2,
32'h1e7de5df,
32'hc6250a18,
32'h584f7b58,
32'hc9edeb50,
32'hc850cab4,
32'hf82a6c6a,
32'h1a4608ab,
32'hc78e9a1d,
32'h57cc15bc,
32'hc91af976,
32'hc337a8f7,
32'hfcdc1342,
32'h15fdf758,
32'hc91af976,
32'h573b2635,
32'hc8507ea7,
32'hbe72d9df,
32'h0192155f,
32'h11a855df,
32'hcac933ae,
32'h569cc31b,
32'hc78e9a1d,
32'hba08fb09,
32'h0645e9af,
32'h0d47d096,
32'hcc983f70,
32'h55f104dc,
32'hc6d569be,
32'hb6002be9,
32'h0af10a22,
32'h08df1a8c,
32'hce86ff2a,
32'h553805f2,
32'hc6250a18,
32'hb25e054b,
32'h0f8cfcbe,
32'h0470ebdc,
32'hd09441bb,
32'h5471e2e6,
32'hc57d965d,
32'haf279193,
32'h14135c94,
32'h00000000,
32'hd2bec333,
32'h539eba45,
32'hc4df2862,
32'hac6145bb,
32'h187de2a7,
32'hfb8f1424,
32'hd5052d97,
32'h52beac9f,
32'hc449d892,
32'haa0efb24,
32'h1cc66e99,
32'hf720e574,
32'hd76619b6,
32'h51d1dc80,
32'hc3bdbdf6,
32'ha833ea44,
32'h20e70f32,
32'hf2b82f6a,
32'hd9e01006,
32'h50d86e6d,
32'hc33aee27,
32'ha6d2a626,
32'h24da0a9a,
32'hee57aa21,
32'hdc71898d,
32'h4fd288dc,
32'hc2c17d52,
32'ha5ed18e0,
32'h2899e64a,
32'hea0208a8,
32'hdf18f0ce,
32'h4ec05432,
32'hc2517e31,
32'ha58480e6,
32'h2c216eaa,
32'he5b9f755,
32'he1d4a2c8,
32'h4da1fab5,
32'hc1eb0209,
32'ha5996f52,
32'h2f6bbe45,
32'he1821a21,
32'he4a2eff6,
32'h4c77a88e,
32'hc18e18a7,
32'ha62bc71b,
32'h32744493,
32'hdd5d0b08,
32'he7821d59,
32'h4b418bbe,
32'hc13ad060,
32'ha73abd3b,
32'h3536cc52,
32'hd94d586c,
32'hea70658a,
32'h49ffd417,
32'hc0f1360b,
32'ha8c4d9cb,
32'h37af8159,
32'hd5558381,
32'hed6bf9d1,
32'h48b2b335,
32'hc0b15502,
32'haac7fa0e,
32'h39daf5e8,
32'hd177fec6,
32'hf0730342,
32'h475a5c77,
32'hc07b371e,
32'had415361,
32'h3bb6276e,
32'hcdb72c7e,
32'hf383a3e2,
32'h45f704f7,
32'hc04ee4b8,
32'hb02d7724,
32'h3d3e82ae,
32'hca155d39,
32'hf69bf7c9,
32'h4488e37f,
32'hc02c64a6,
32'hb3885772,
32'h3e71e759,
32'hc694ce67,
32'hf9ba1651,
32'h43103085,
32'hc013bc39,
32'hb74d4ccb,
32'h3f4eaafe,
32'hc337a8f7,
32'hfcdc1342,
32'h418d2621,
32'hc004ef3f,
32'hbb771c81,
32'h3fd39b5a
};

always @(posedge clk) 
  if (en)
    dout <= mem[addr];

endmodule

/*
const int twidTabEven[4*6 + 16*6 + 64*6] = {
	0x40000000, 0x00000000, 0x40000000, 0x00000000, 0x40000000, 0x00000000, 0x5a82799a, 0xd2bec333, 
	0x539eba45, 0xe7821d59, 0x539eba45, 0xc4df2862, 0x40000000, 0xc0000000, 0x5a82799a, 0xd2bec333, 
	0x00000000, 0xd2bec333, 0x00000000, 0xd2bec333, 0x539eba45, 0xc4df2862, 0xac6145bb, 0x187de2a7, 
	
	0x40000000, 0x00000000, 0x40000000, 0x00000000, 0x40000000, 0x00000000, 0x4b418bbe, 0xf383a3e2, 
	0x45f704f7, 0xf9ba1651, 0x4fd288dc, 0xed6bf9d1, 0x539eba45, 0xe7821d59, 0x4b418bbe, 0xf383a3e2, 
	0x58c542c5, 0xdc71898d, 0x58c542c5, 0xdc71898d, 0x4fd288dc, 0xed6bf9d1, 0x5a12e720, 0xce86ff2a, 
	0x5a82799a, 0xd2bec333, 0x539eba45, 0xe7821d59, 0x539eba45, 0xc4df2862, 0x58c542c5, 0xcac933ae, 
	0x569cc31b, 0xe1d4a2c8, 0x45f704f7, 0xc04ee4b8, 0x539eba45, 0xc4df2862, 0x58c542c5, 0xdc71898d, 
	0x3248d382, 0xc13ad060, 0x4b418bbe, 0xc13ad060, 0x5a12e720, 0xd76619b6, 0x1a4608ab, 0xc78e9a1d, 
	0x40000000, 0xc0000000, 0x5a82799a, 0xd2bec333, 0x00000000, 0xd2bec333, 0x3248d382, 0xc13ad060, 
	0x5a12e720, 0xce86ff2a, 0xe5b9f755, 0xe1d4a2c8, 0x22a2f4f8, 0xc4df2862, 0x58c542c5, 0xcac933ae, 
	0xcdb72c7e, 0xf383a3e2, 0x11a855df, 0xcac933ae, 0x569cc31b, 0xc78e9a1d, 0xba08fb09, 0x0645e9af, 
	0x00000000, 0xd2bec333, 0x539eba45, 0xc4df2862, 0xac6145bb, 0x187de2a7, 0xee57aa21, 0xdc71898d, 
	0x4fd288dc, 0xc2c17d52, 0xa5ed18e0, 0x2899e64a, 0xdd5d0b08, 0xe7821d59, 0x4b418bbe, 0xc13ad060, 
	0xa73abd3b, 0x3536cc52, 0xcdb72c7e, 0xf383a3e2, 0x45f704f7, 0xc04ee4b8, 0xb02d7724, 0x3d3e82ae, 
	
	0x40000000, 0x00000000, 0x40000000, 0x00000000, 0x40000000, 0x00000000, 0x43103085, 0xfcdc1342, 
	0x418d2621, 0xfe6deaa1, 0x4488e37f, 0xfb4ab7db, 0x45f704f7, 0xf9ba1651, 0x43103085, 0xfcdc1342, 
	0x48b2b335, 0xf69bf7c9, 0x48b2b335, 0xf69bf7c9, 0x4488e37f, 0xfb4ab7db, 0x4c77a88e, 0xf1fa3ecb, 
	0x4b418bbe, 0xf383a3e2, 0x45f704f7, 0xf9ba1651, 0x4fd288dc, 0xed6bf9d1, 0x4da1fab5, 0xf0730342, 
	0x475a5c77, 0xf82a6c6a, 0x52beac9f, 0xe8f77acf, 0x4fd288dc, 0xed6bf9d1, 0x48b2b335, 0xf69bf7c9, 
	0x553805f2, 0xe4a2eff6, 0x51d1dc80, 0xea70658a, 0x49ffd417, 0xf50ef5de, 0x573b2635, 0xe0745b24, 
	0x539eba45, 0xe7821d59, 0x4b418bbe, 0xf383a3e2, 0x58c542c5, 0xdc71898d, 0x553805f2, 0xe4a2eff6, 
	0x4c77a88e, 0xf1fa3ecb, 0x59d438e5, 0xd8a00bae, 0x569cc31b, 0xe1d4a2c8, 0x4da1fab5, 0xf0730342, 
	0x5a6690ae, 0xd5052d97, 0x57cc15bc, 0xdf18f0ce, 0x4ec05432, 0xeeee2d9d, 0x5a7b7f1a, 0xd1a5ef90, 
	0x58c542c5, 0xdc71898d, 0x4fd288dc, 0xed6bf9d1, 0x5a12e720, 0xce86ff2a, 0x5987b08a, 0xd9e01006, 
	0x50d86e6d, 0xebeca36c, 0x592d59da, 0xcbacb0bf, 0x5a12e720, 0xd76619b6, 0x51d1dc80, 0xea70658a, 
	0x57cc15bc, 0xc91af976, 0x5a6690ae, 0xd5052d97, 0x52beac9f, 0xe8f77acf, 0x55f104dc, 0xc6d569be, 
	0x5a82799a, 0xd2bec333, 0x539eba45, 0xe7821d59, 0x539eba45, 0xc4df2862, 0x5a6690ae, 0xd09441bb, 
	0x5471e2e6, 0xe61086bc, 0x50d86e6d, 0xc33aee27, 0x5a12e720, 0xce86ff2a, 0x553805f2, 0xe4a2eff6, 
	0x4da1fab5, 0xc1eb0209, 0x5987b08a, 0xcc983f70, 0x55f104dc, 0xe3399167, 0x49ffd417, 0xc0f1360b, 
	0x58c542c5, 0xcac933ae, 0x569cc31b, 0xe1d4a2c8, 0x45f704f7, 0xc04ee4b8, 0x57cc15bc, 0xc91af976, 
	0x573b2635, 0xe0745b24, 0x418d2621, 0xc004ef3f, 0x569cc31b, 0xc78e9a1d, 0x57cc15bc, 0xdf18f0ce, 
	0x3cc85709, 0xc013bc39, 0x553805f2, 0xc6250a18, 0x584f7b58, 0xddc29958, 0x37af354c, 0xc07b371e, 
	0x539eba45, 0xc4df2862, 0x58c542c5, 0xdc71898d, 0x3248d382, 0xc13ad060, 0x51d1dc80, 0xc3bdbdf6, 
	0x592d59da, 0xdb25f566, 0x2c9caf6c, 0xc2517e31, 0x4fd288dc, 0xc2c17d52, 0x5987b08a, 0xd9e01006, 
	0x26b2a794, 0xc3bdbdf6, 0x4da1fab5, 0xc1eb0209, 0x59d438e5, 0xd8a00bae, 0x2092f05f, 0xc57d965d, 
	0x4b418bbe, 0xc13ad060, 0x5a12e720, 0xd76619b6, 0x1a4608ab, 0xc78e9a1d, 0x48b2b335, 0xc0b15502, 
	0x5a43b190, 0xd6326a88, 0x13d4ae08, 0xc9edeb50, 0x45f704f7, 0xc04ee4b8, 0x5a6690ae, 0xd5052d97, 
	0x0d47d096, 0xcc983f70, 0x43103085, 0xc013bc39, 0x5a7b7f1a, 0xd3de9156, 0x06a886a0, 0xcf89e3e8, 
	0x40000000, 0xc0000000, 0x5a82799a, 0xd2bec333, 0x00000000, 0xd2bec333, 0x3cc85709, 0xc013bc39, 
	0x5a7b7f1a, 0xd1a5ef90, 0xf9577960, 0xd6326a88, 0x396b3199, 0xc04ee4b8, 0x5a6690ae, 0xd09441bb, 
	0xf2b82f6a, 0xd9e01006, 0x35eaa2c7, 0xc0b15502, 0x5a43b190, 0xcf89e3e8, 0xec2b51f8, 0xddc29958, 
	0x3248d382, 0xc13ad060, 0x5a12e720, 0xce86ff2a, 0xe5b9f755, 0xe1d4a2c8, 0x2e88013a, 0xc1eb0209, 
	0x59d438e5, 0xcd8bbb6d, 0xdf6d0fa1, 0xe61086bc, 0x2aaa7c7f, 0xc2c17d52, 0x5987b08a, 0xcc983f70, 
	0xd94d586c, 0xea70658a, 0x26b2a794, 0xc3bdbdf6, 0x592d59da, 0xcbacb0bf, 0xd3635094, 0xeeee2d9d, 
	0x22a2f4f8, 0xc4df2862, 0x58c542c5, 0xcac933ae, 0xcdb72c7e, 0xf383a3e2, 0x1e7de5df, 0xc6250a18, 
	0x584f7b58, 0xc9edeb50, 0xc850cab4, 0xf82a6c6a, 0x1a4608ab, 0xc78e9a1d, 0x57cc15bc, 0xc91af976, 
	0xc337a8f7, 0xfcdc1342, 0x15fdf758, 0xc91af976, 0x573b2635, 0xc8507ea7, 0xbe72d9df, 0x0192155f, 
	0x11a855df, 0xcac933ae, 0x569cc31b, 0xc78e9a1d, 0xba08fb09, 0x0645e9af, 0x0d47d096, 0xcc983f70, 
	0x55f104dc, 0xc6d569be, 0xb6002be9, 0x0af10a22, 0x08df1a8c, 0xce86ff2a, 0x553805f2, 0xc6250a18, 
	0xb25e054b, 0x0f8cfcbe, 0x0470ebdc, 0xd09441bb, 0x5471e2e6, 0xc57d965d, 0xaf279193, 0x14135c94, 
	0x00000000, 0xd2bec333, 0x539eba45, 0xc4df2862, 0xac6145bb, 0x187de2a7, 0xfb8f1424, 0xd5052d97, 
	0x52beac9f, 0xc449d892, 0xaa0efb24, 0x1cc66e99, 0xf720e574, 0xd76619b6, 0x51d1dc80, 0xc3bdbdf6, 
	0xa833ea44, 0x20e70f32, 0xf2b82f6a, 0xd9e01006, 0x50d86e6d, 0xc33aee27, 0xa6d2a626, 0x24da0a9a, 
	0xee57aa21, 0xdc71898d, 0x4fd288dc, 0xc2c17d52, 0xa5ed18e0, 0x2899e64a, 0xea0208a8, 0xdf18f0ce, 
	0x4ec05432, 0xc2517e31, 0xa58480e6, 0x2c216eaa, 0xe5b9f755, 0xe1d4a2c8, 0x4da1fab5, 0xc1eb0209, 
	0xa5996f52, 0x2f6bbe45, 0xe1821a21, 0xe4a2eff6, 0x4c77a88e, 0xc18e18a7, 0xa62bc71b, 0x32744493, 
	0xdd5d0b08, 0xe7821d59, 0x4b418bbe, 0xc13ad060, 0xa73abd3b, 0x3536cc52, 0xd94d586c, 0xea70658a, 
	0x49ffd417, 0xc0f1360b, 0xa8c4d9cb, 0x37af8159, 0xd5558381, 0xed6bf9d1, 0x48b2b335, 0xc0b15502, 
	0xaac7fa0e, 0x39daf5e8, 0xd177fec6, 0xf0730342, 0x475a5c77, 0xc07b371e, 0xad415361, 0x3bb6276e, 
	0xcdb72c7e, 0xf383a3e2, 0x45f704f7, 0xc04ee4b8, 0xb02d7724, 0x3d3e82ae, 0xca155d39, 0xf69bf7c9, 
	0x4488e37f, 0xc02c64a6, 0xb3885772, 0x3e71e759, 0xc694ce67, 0xf9ba1651, 0x43103085, 0xc013bc39, 
	0xb74d4ccb, 0x3f4eaafe, 0xc337a8f7, 0xfcdc1342, 0x418d2621, 0xc004ef3f, 0xbb771c81, 0x3fd39b5a, 
};


*/
