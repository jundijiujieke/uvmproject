module rom_twidTabOdd(
clk,
en,
addr,

dout
);

input clk;
input en;
input [9:0] addr;

output reg [31:0] dout;

reg [31:0] mem[0:1009]={ 

32'h40000000,
32'h00000000,
32'h40000000,
32'h00000000,
32'h40000000,
32'h00000000,
32'h539eba45,
32'he7821d59,
32'h4b418bbe,
32'hf383a3e2,
32'h58c542c5,
32'hdc71898d,
32'h5a82799a,
32'hd2bec333,
32'h539eba45,
32'he7821d59,
32'h539eba45,
32'hc4df2862,
32'h539eba45,
32'hc4df2862,
32'h58c542c5,
32'hdc71898d,
32'h3248d382,
32'hc13ad060,
32'h40000000,
32'hc0000000,
32'h5a82799a,
32'hd2bec333,
32'h00000000,
32'hd2bec333,
32'h22a2f4f8,
32'hc4df2862,
32'h58c542c5,
32'hcac933ae,
32'hcdb72c7e,
32'hf383a3e2,
32'h00000000,
32'hd2bec333,
32'h539eba45,
32'hc4df2862,
32'hac6145bb,
32'h187de2a7,
32'hdd5d0b08,
32'he7821d59,
32'h4b418bbe,
32'hc13ad060,
32'ha73abd3b,
32'h3536cc52,
32'h40000000,
32'h00000000,
32'h40000000,
32'h00000000,
32'h40000000,
32'h00000000,
32'h45f704f7,
32'hf9ba1651,
32'h43103085,
32'hfcdc1342,
32'h48b2b335,
32'hf69bf7c9,
32'h4b418bbe,
32'hf383a3e2,
32'h45f704f7,
32'hf9ba1651,
32'h4fd288dc,
32'hed6bf9d1,
32'h4fd288dc,
32'hed6bf9d1,
32'h48b2b335,
32'hf69bf7c9,
32'h553805f2,
32'he4a2eff6,
32'h539eba45,
32'he7821d59,
32'h4b418bbe,
32'hf383a3e2,
32'h58c542c5,
32'hdc71898d,
32'h569cc31b,
32'he1d4a2c8,
32'h4da1fab5,
32'hf0730342,
32'h5a6690ae,
32'hd5052d97,
32'h58c542c5,
32'hdc71898d,
32'h4fd288dc,
32'hed6bf9d1,
32'h5a12e720,
32'hce86ff2a,
32'h5a12e720,
32'hd76619b6,
32'h51d1dc80,
32'hea70658a,
32'h57cc15bc,
32'hc91af976,
32'h5a82799a,
32'hd2bec333,
32'h539eba45,
32'he7821d59,
32'h539eba45,
32'hc4df2862,
32'h5a12e720,
32'hce86ff2a,
32'h553805f2,
32'he4a2eff6,
32'h4da1fab5,
32'hc1eb0209,
32'h58c542c5,
32'hcac933ae,
32'h569cc31b,
32'he1d4a2c8,
32'h45f704f7,
32'hc04ee4b8,
32'h569cc31b,
32'hc78e9a1d,
32'h57cc15bc,
32'hdf18f0ce,
32'h3cc85709,
32'hc013bc39,
32'h539eba45,
32'hc4df2862,
32'h58c542c5,
32'hdc71898d,
32'h3248d382,
32'hc13ad060,
32'h4fd288dc,
32'hc2c17d52,
32'h5987b08a,
32'hd9e01006,
32'h26b2a794,
32'hc3bdbdf6,
32'h4b418bbe,
32'hc13ad060,
32'h5a12e720,
32'hd76619b6,
32'h1a4608ab,
32'hc78e9a1d,
32'h45f704f7,
32'hc04ee4b8,
32'h5a6690ae,
32'hd5052d97,
32'h0d47d096,
32'hcc983f70,
32'h40000000,
32'hc0000000,
32'h5a82799a,
32'hd2bec333,
32'h00000000,
32'hd2bec333,
32'h396b3199,
32'hc04ee4b8,
32'h5a6690ae,
32'hd09441bb,
32'hf2b82f6a,
32'hd9e01006,
32'h3248d382,
32'hc13ad060,
32'h5a12e720,
32'hce86ff2a,
32'he5b9f755,
32'he1d4a2c8,
32'h2aaa7c7f,
32'hc2c17d52,
32'h5987b08a,
32'hcc983f70,
32'hd94d586c,
32'hea70658a,
32'h22a2f4f8,
32'hc4df2862,
32'h58c542c5,
32'hcac933ae,
32'hcdb72c7e,
32'hf383a3e2,
32'h1a4608ab,
32'hc78e9a1d,
32'h57cc15bc,
32'hc91af976,
32'hc337a8f7,
32'hfcdc1342,
32'h11a855df,
32'hcac933ae,
32'h569cc31b,
32'hc78e9a1d,
32'hba08fb09,
32'h0645e9af,
32'h08df1a8c,
32'hce86ff2a,
32'h553805f2,
32'hc6250a18,
32'hb25e054b,
32'h0f8cfcbe,
32'h00000000,
32'hd2bec333,
32'h539eba45,
32'hc4df2862,
32'hac6145bb,
32'h187de2a7,
32'hf720e574,
32'hd76619b6,
32'h51d1dc80,
32'hc3bdbdf6,
32'ha833ea44,
32'h20e70f32,
32'hee57aa21,
32'hdc71898d,
32'h4fd288dc,
32'hc2c17d52,
32'ha5ed18e0,
32'h2899e64a,
32'he5b9f755,
32'he1d4a2c8,
32'h4da1fab5,
32'hc1eb0209,
32'ha5996f52,
32'h2f6bbe45,
32'hdd5d0b08,
32'he7821d59,
32'h4b418bbe,
32'hc13ad060,
32'ha73abd3b,
32'h3536cc52,
32'hd5558381,
32'hed6bf9d1,
32'h48b2b335,
32'hc0b15502,
32'haac7fa0e,
32'h39daf5e8,
32'hcdb72c7e,
32'hf383a3e2,
32'h45f704f7,
32'hc04ee4b8,
32'hb02d7724,
32'h3d3e82ae,
32'hc694ce67,
32'hf9ba1651,
32'h43103085,
32'hc013bc39,
32'hb74d4ccb,
32'h3f4eaafe,
32'h40000000,
32'h00000000,
32'h40000000,
32'h00000000,
32'h40000000,
32'h00000000,
32'h418d2621,
32'hfe6deaa1,
32'h40c7d2bd,
32'hff36f170,
32'h424ff28f,
32'hfda4f351,
32'h43103085,
32'hfcdc1342,
32'h418d2621,
32'hfe6deaa1,
32'h4488e37f,
32'hfb4ab7db,
32'h4488e37f,
32'hfb4ab7db,
32'h424ff28f,
32'hfda4f351,
32'h46aa0d6d,
32'hf8f21e8e,
32'h45f704f7,
32'hf9ba1651,
32'h43103085,
32'hfcdc1342,
32'h48b2b335,
32'hf69bf7c9,
32'h475a5c77,
32'hf82a6c6a,
32'h43cdd89a,
32'hfc135231,
32'h4aa22036,
32'hf4491311,
32'h48b2b335,
32'hf69bf7c9,
32'h4488e37f,
32'hfb4ab7db,
32'h4c77a88e,
32'hf1fa3ecb,
32'h49ffd417,
32'hf50ef5de,
32'h454149fc,
32'hfa824bfd,
32'h4e32a956,
32'hefb047f2,
32'h4b418bbe,
32'hf383a3e2,
32'h45f704f7,
32'hf9ba1651,
32'h4fd288dc,
32'hed6bf9d1,
32'h4c77a88e,
32'hf1fa3ecb,
32'h46aa0d6d,
32'hf8f21e8e,
32'h5156b6d9,
32'heb2e1dbe,
32'h4da1fab5,
32'hf0730342,
32'h475a5c77,
32'hf82a6c6a,
32'h52beac9f,
32'he8f77acf,
32'h4ec05432,
32'heeee2d9d,
32'h4807eb4b,
32'hf7630799,
32'h5409ed4b,
32'he6c8d59c,
32'h4fd288dc,
32'hed6bf9d1,
32'h48b2b335,
32'hf69bf7c9,
32'h553805f2,
32'he4a2eff6,
32'h50d86e6d,
32'hebeca36c,
32'h495aada2,
32'hf5d544a7,
32'h56488dc5,
32'he28688a4,
32'h51d1dc80,
32'hea70658a,
32'h49ffd417,
32'hf50ef5de,
32'h573b2635,
32'he0745b24,
32'h52beac9f,
32'he8f77acf,
32'h4aa22036,
32'hf4491311,
32'h580f7b19,
32'hde6d1f65,
32'h539eba45,
32'he7821d59,
32'h4b418bbe,
32'hf383a3e2,
32'h58c542c5,
32'hdc71898d,
32'h5471e2e6,
32'he61086bc,
32'h4bde1089,
32'hf2beafed,
32'h595c3e2a,
32'hda8249b4,
32'h553805f2,
32'he4a2eff6,
32'h4c77a88e,
32'hf1fa3ecb,
32'h59d438e5,
32'hd8a00bae,
32'h55f104dc,
32'he3399167,
32'h4d0e4de2,
32'hf136580d,
32'h5a2d0957,
32'hd6cb76c9,
32'h569cc31b,
32'he1d4a2c8,
32'h4da1fab5,
32'hf0730342,
32'h5a6690ae,
32'hd5052d97,
32'h573b2635,
32'he0745b24,
32'h4e32a956,
32'hefb047f2,
32'h5a80baf6,
32'hd34dcdb4,
32'h57cc15bc,
32'hdf18f0ce,
32'h4ec05432,
32'heeee2d9d,
32'h5a7b7f1a,
32'hd1a5ef90,
32'h584f7b58,
32'hddc29958,
32'h4f4af5d1,
32'hee2cbbc1,
32'h5a56deec,
32'hd00e2639,
32'h58c542c5,
32'hdc71898d,
32'h4fd288dc,
32'hed6bf9d1,
32'h5a12e720,
32'hce86ff2a,
32'h592d59da,
32'hdb25f566,
32'h50570819,
32'hecabef3d,
32'h59afaf4c,
32'hcd110216,
32'h5987b08a,
32'hd9e01006,
32'h50d86e6d,
32'hebeca36c,
32'h592d59da,
32'hcbacb0bf,
32'h59d438e5,
32'hd8a00bae,
32'h5156b6d9,
32'heb2e1dbe,
32'h588c1404,
32'hca5a86c4,
32'h5a12e720,
32'hd76619b6,
32'h51d1dc80,
32'hea70658a,
32'h57cc15bc,
32'hc91af976,
32'h5a43b190,
32'hd6326a88,
32'h5249daa2,
32'he9b38223,
32'h56eda1a0,
32'hc7ee77b3,
32'h5a6690ae,
32'hd5052d97,
32'h52beac9f,
32'he8f77acf,
32'h55f104dc,
32'hc6d569be,
32'h5a7b7f1a,
32'hd3de9156,
32'h53304df6,
32'he83c56cf,
32'h54d69714,
32'hc5d03118,
32'h5a82799a,
32'hd2bec333,
32'h539eba45,
32'he7821d59,
32'h539eba45,
32'hc4df2862,
32'h5a7b7f1a,
32'hd1a5ef90,
32'h5409ed4b,
32'he6c8d59c,
32'h5249daa2,
32'hc402a33c,
32'h5a6690ae,
32'hd09441bb,
32'h5471e2e6,
32'he61086bc,
32'h50d86e6d,
32'hc33aee27,
32'h5a43b190,
32'hcf89e3e8,
32'h54d69714,
32'he55937d5,
32'h4f4af5d1,
32'hc2884e6e,
32'h5a12e720,
32'hce86ff2a,
32'h553805f2,
32'he4a2eff6,
32'h4da1fab5,
32'hc1eb0209,
32'h59d438e5,
32'hcd8bbb6d,
32'h55962bc0,
32'he3edb628,
32'h4bde1089,
32'hc1633f8a,
32'h5987b08a,
32'hcc983f70,
32'h55f104dc,
32'he3399167,
32'h49ffd417,
32'hc0f1360b,
32'h592d59da,
32'hcbacb0bf,
32'h56488dc5,
32'he28688a4,
32'h4807eb4b,
32'hc0950d1d,
32'h58c542c5,
32'hcac933ae,
32'h569cc31b,
32'he1d4a2c8,
32'h45f704f7,
32'hc04ee4b8,
32'h584f7b58,
32'hc9edeb50,
32'h56eda1a0,
32'he123e6ad,
32'h43cdd89a,
32'hc01ed535,
32'h57cc15bc,
32'hc91af976,
32'h573b2635,
32'he0745b24,
32'h418d2621,
32'hc004ef3f,
32'h573b2635,
32'hc8507ea7,
32'h57854ddd,
32'hdfc606f1,
32'h3f35b59d,
32'hc0013bd3,
32'h569cc31b,
32'hc78e9a1d,
32'h57cc15bc,
32'hdf18f0ce,
32'h3cc85709,
32'hc013bc39,
32'h55f104dc,
32'hc6d569be,
32'h580f7b19,
32'hde6d1f65,
32'h3a45e1f7,
32'hc03c6a07,
32'h553805f2,
32'hc6250a18,
32'h584f7b58,
32'hddc29958,
32'h37af354c,
32'hc07b371e,
32'h5471e2e6,
32'hc57d965d,
32'h588c1404,
32'hdd196538,
32'h350536f1,
32'hc0d00db6,
32'h539eba45,
32'hc4df2862,
32'h58c542c5,
32'hdc71898d,
32'h3248d382,
32'hc13ad060,
32'h52beac9f,
32'hc449d892,
32'h58fb0568,
32'hdbcb0cce,
32'h2f7afdfc,
32'hc1bb5a11,
32'h51d1dc80,
32'hc3bdbdf6,
32'h592d59da,
32'hdb25f566,
32'h2c9caf6c,
32'hc2517e31,
32'h50d86e6d,
32'hc33aee27,
32'h595c3e2a,
32'hda8249b4,
32'h29aee694,
32'hc2fd08a9,
32'h4fd288dc,
32'hc2c17d52,
32'h5987b08a,
32'hd9e01006,
32'h26b2a794,
32'hc3bdbdf6,
32'h4ec05432,
32'hc2517e31,
32'h59afaf4c,
32'hd93f4e9e,
32'h23a8fb93,
32'hc4935b3c,
32'h4da1fab5,
32'hc1eb0209,
32'h59d438e5,
32'hd8a00bae,
32'h2092f05f,
32'hc57d965d,
32'h4c77a88e,
32'hc18e18a7,
32'h59f54bee,
32'hd8024d59,
32'h1d719810,
32'hc67c1e18,
32'h4b418bbe,
32'hc13ad060,
32'h5a12e720,
32'hd76619b6,
32'h1a4608ab,
32'hc78e9a1d,
32'h49ffd417,
32'hc0f1360b,
32'h5a2d0957,
32'hd6cb76c9,
32'h17115bc0,
32'hc8b4ab32,
32'h48b2b335,
32'hc0b15502,
32'h5a43b190,
32'hd6326a88,
32'h13d4ae08,
32'hc9edeb50,
32'h475a5c77,
32'hc07b371e,
32'h5a56deec,
32'hd59afadb,
32'h10911f04,
32'hcb39edca,
32'h45f704f7,
32'hc04ee4b8,
32'h5a6690ae,
32'hd5052d97,
32'h0d47d096,
32'hcc983f70,
32'h4488e37f,
32'hc02c64a6,
32'h5a72c63b,
32'hd4710883,
32'h09f9e6a1,
32'hce0866b8,
32'h43103085,
32'hc013bc39,
32'h5a7b7f1a,
32'hd3de9156,
32'h06a886a0,
32'hcf89e3e8,
32'h418d2621,
32'hc004ef3f,
32'h5a80baf6,
32'hd34dcdb4,
32'h0354d741,
32'hd11c3142,
32'h40000000,
32'hc0000000,
32'h5a82799a,
32'hd2bec333,
32'h00000000,
32'hd2bec333,
32'h3e68fb62,
32'hc004ef3f,
32'h5a80baf6,
32'hd2317756,
32'hfcab28bf,
32'hd4710883,
32'h3cc85709,
32'hc013bc39,
32'h5a7b7f1a,
32'hd1a5ef90,
32'hf9577960,
32'hd6326a88,
32'h3b1e5335,
32'hc02c64a6,
32'h5a72c63b,
32'hd11c3142,
32'hf606195f,
32'hd8024d59,
32'h396b3199,
32'hc04ee4b8,
32'h5a6690ae,
32'hd09441bb,
32'hf2b82f6a,
32'hd9e01006,
32'h37af354c,
32'hc07b371e,
32'h5a56deec,
32'hd00e2639,
32'hef6ee0fc,
32'hdbcb0cce,
32'h35eaa2c7,
32'hc0b15502,
32'h5a43b190,
32'hcf89e3e8,
32'hec2b51f8,
32'hddc29958,
32'h341dbfd3,
32'hc0f1360b,
32'h5a2d0957,
32'hcf077fe1,
32'he8eea440,
32'hdfc606f1,
32'h3248d382,
32'hc13ad060,
32'h5a12e720,
32'hce86ff2a,
32'he5b9f755,
32'he1d4a2c8,
32'h306c2624,
32'hc18e18a7,
32'h59f54bee,
32'hce0866b8,
32'he28e67f0,
32'he3edb628,
32'h2e88013a,
32'hc1eb0209,
32'h59d438e5,
32'hcd8bbb6d,
32'hdf6d0fa1,
32'he61086bc,
32'h2c9caf6c,
32'hc2517e31,
32'h59afaf4c,
32'hcd110216,
32'hdc57046d,
32'he83c56cf,
32'h2aaa7c7f,
32'hc2c17d52,
32'h5987b08a,
32'hcc983f70,
32'hd94d586c,
32'hea70658a,
32'h28b1b544,
32'hc33aee27,
32'h595c3e2a,
32'hcc217822,
32'hd651196c,
32'hecabef3d,
32'h26b2a794,
32'hc3bdbdf6,
32'h592d59da,
32'hcbacb0bf,
32'hd3635094,
32'heeee2d9d,
32'h24ada23d,
32'hc449d892,
32'h58fb0568,
32'hcb39edca,
32'hd0850204,
32'hf136580d,
32'h22a2f4f8,
32'hc4df2862,
32'h58c542c5,
32'hcac933ae,
32'hcdb72c7e,
32'hf383a3e2,
32'h2092f05f,
32'hc57d965d,
32'h588c1404,
32'hca5a86c4,
32'hcafac90f,
32'hf5d544a7,
32'h1e7de5df,
32'hc6250a18,
32'h584f7b58,
32'hc9edeb50,
32'hc850cab4,
32'hf82a6c6a,
32'h1c6427a9,
32'hc6d569be,
32'h580f7b19,
32'hc9836582,
32'hc5ba1e09,
32'hfa824bfd,
32'h1a4608ab,
32'hc78e9a1d,
32'h57cc15bc,
32'hc91af976,
32'hc337a8f7,
32'hfcdc1342,
32'h1823dc7d,
32'hc8507ea7,
32'h57854ddd,
32'hc8b4ab32,
32'hc0ca4a63,
32'hff36f170,
32'h15fdf758,
32'hc91af976,
32'h573b2635,
32'hc8507ea7,
32'hbe72d9df,
32'h0192155f,
32'h13d4ae08,
32'hc9edeb50,
32'h56eda1a0,
32'hc7ee77b3,
32'hbc322766,
32'h03ecadcf,
32'h11a855df,
32'hcac933ae,
32'h569cc31b,
32'hc78e9a1d,
32'hba08fb09,
32'h0645e9af,
32'h0f7944a7,
32'hcbacb0bf,
32'h56488dc5,
32'hc730e997,
32'hb7f814b5,
32'h089cf867,
32'h0d47d096,
32'hcc983f70,
32'h55f104dc,
32'hc6d569be,
32'hb6002be9,
32'h0af10a22,
32'h0b145041,
32'hcd8bbb6d,
32'h55962bc0,
32'hc67c1e18,
32'hb421ef77,
32'h0d415013,
32'h08df1a8c,
32'hce86ff2a,
32'h553805f2,
32'hc6250a18,
32'hb25e054b,
32'h0f8cfcbe,
32'h06a886a0,
32'hcf89e3e8,
32'h54d69714,
32'hc5d03118,
32'hb0b50a2f,
32'h11d3443f,
32'h0470ebdc,
32'hd09441bb,
32'h5471e2e6,
32'hc57d965d,
32'haf279193,
32'h14135c94,
32'h0238a1c6,
32'hd1a5ef90,
32'h5409ed4b,
32'hc52d3d18,
32'hadb6255e,
32'h164c7ddd,
32'h00000000,
32'hd2bec333,
32'h539eba45,
32'hc4df2862,
32'hac6145bb,
32'h187de2a7,
32'hfdc75e3a,
32'hd3de9156,
32'h53304df6,
32'hc4935b3c,
32'hab2968ec,
32'h1aa6c82b,
32'hfb8f1424,
32'hd5052d97,
32'h52beac9f,
32'hc449d892,
32'haa0efb24,
32'h1cc66e99,
32'hf9577960,
32'hd6326a88,
32'h5249daa2,
32'hc402a33c,
32'ha9125e60,
32'h1edc1953,
32'hf720e574,
32'hd76619b6,
32'h51d1dc80,
32'hc3bdbdf6,
32'ha833ea44,
32'h20e70f32,
32'hf4ebafbf,
32'hd8a00bae,
32'h5156b6d9,
32'hc37b2b6a,
32'ha773ebfc,
32'h22e69ac8,
32'hf2b82f6a,
32'hd9e01006,
32'h50d86e6d,
32'hc33aee27,
32'ha6d2a626,
32'h24da0a9a,
32'hf086bb59,
32'hdb25f566,
32'h50570819,
32'hc2fd08a9,
32'ha65050b4,
32'h26c0b162,
32'hee57aa21,
32'hdc71898d,
32'h4fd288dc,
32'hc2c17d52,
32'ha5ed18e0,
32'h2899e64a,
32'hec2b51f8,
32'hddc29958,
32'h4f4af5d1,
32'hc2884e6e,
32'ha5a92114,
32'h2a650525,
32'hea0208a8,
32'hdf18f0ce,
32'h4ec05432,
32'hc2517e31,
32'ha58480e6,
32'h2c216eaa,
32'he7dc2383,
32'he0745b24,
32'h4e32a956,
32'hc21d0eb8,
32'ha57f450a,
32'h2dce88aa,
32'he5b9f755,
32'he1d4a2c8,
32'h4da1fab5,
32'hc1eb0209,
32'ha5996f52,
32'h2f6bbe45,
32'he39bd857,
32'he3399167,
32'h4d0e4de2,
32'hc1bb5a11,
32'ha5d2f6a9,
32'h30f8801f,
32'he1821a21,
32'he4a2eff6,
32'h4c77a88e,
32'hc18e18a7,
32'ha62bc71b,
32'h32744493,
32'hdf6d0fa1,
32'he61086bc,
32'h4bde1089,
32'hc1633f8a,
32'ha6a3c1d6,
32'h33de87de,
32'hdd5d0b08,
32'he7821d59,
32'h4b418bbe,
32'hc13ad060,
32'ha73abd3b,
32'h3536cc52,
32'hdb525dc3,
32'he8f77acf,
32'h4aa22036,
32'hc114ccb9,
32'ha7f084e7,
32'h367c9a7e,
32'hd94d586c,
32'hea70658a,
32'h49ffd417,
32'hc0f1360b,
32'ha8c4d9cb,
32'h37af8159,
32'hd74e4abc,
32'hebeca36c,
32'h495aada2,
32'hc0d00db6,
32'ha9b7723b,
32'h38cf1669,
32'hd5558381,
32'hed6bf9d1,
32'h48b2b335,
32'hc0b15502,
32'haac7fa0e,
32'h39daf5e8,
32'hd3635094,
32'heeee2d9d,
32'h4807eb4b,
32'hc0950d1d,
32'habf612b5,
32'h3ad2c2e8,
32'hd177fec6,
32'hf0730342,
32'h475a5c77,
32'hc07b371e,
32'had415361,
32'h3bb6276e,
32'hcf93d9dc,
32'hf1fa3ecb,
32'h46aa0d6d,
32'hc063d405,
32'haea94927,
32'h3c84d496,
32'hcdb72c7e,
32'hf383a3e2,
32'h45f704f7,
32'hc04ee4b8,
32'hb02d7724,
32'h3d3e82ae,
32'hcbe2402d,
32'hf50ef5de,
32'h454149fc,
32'hc03c6a07,
32'hb1cd56aa,
32'h3de2f148,
32'hca155d39,
32'hf69bf7c9,
32'h4488e37f,
32'hc02c64a6,
32'hb3885772,
32'h3e71e759,
32'hc850cab4,
32'hf82a6c6a,
32'h43cdd89a,
32'hc01ed535,
32'hb55ddfca,
32'h3eeb3347,
32'hc694ce67,
32'hf9ba1651,
32'h43103085,
32'hc013bc39,
32'hb74d4ccb,
32'h3f4eaafe,
32'hc4e1accb,
32'hfb4ab7db,
32'h424ff28f,
32'hc00b1a20,
32'hb955f293,
32'h3f9c2bfb,
32'hc337a8f7,
32'hfcdc1342,
32'h418d2621,
32'hc004ef3f,
32'hbb771c81,
32'h3fd39b5a,
32'hc197049e,
32'hfe6deaa1,
32'h40c7d2bd,
32'hc0013bd3,
32'hbdb00d71,
32'h3ff4e5e0,
32'h00000000,
32'h00000000
};

always @(posedge clk) 
  if (en)
    dout <= mem[addr];

endmodule
/*
const int twidTabOdd[8*6 + 32*6 + 128*6] = {
	0x40000000, 0x00000000, 0x40000000, 0x00000000, 0x40000000, 0x00000000, 0x539eba45, 0xe7821d59, 
	0x4b418bbe, 0xf383a3e2, 0x58c542c5, 0xdc71898d, 0x5a82799a, 0xd2bec333, 0x539eba45, 0xe7821d59, 
	0x539eba45, 0xc4df2862, 0x539eba45, 0xc4df2862, 0x58c542c5, 0xdc71898d, 0x3248d382, 0xc13ad060, 
	0x40000000, 0xc0000000, 0x5a82799a, 0xd2bec333, 0x00000000, 0xd2bec333, 0x22a2f4f8, 0xc4df2862, 
	0x58c542c5, 0xcac933ae, 0xcdb72c7e, 0xf383a3e2, 0x00000000, 0xd2bec333, 0x539eba45, 0xc4df2862, 
	0xac6145bb, 0x187de2a7, 0xdd5d0b08, 0xe7821d59, 0x4b418bbe, 0xc13ad060, 0xa73abd3b, 0x3536cc52, 
	
	0x40000000, 0x00000000, 0x40000000, 0x00000000, 0x40000000, 0x00000000, 0x45f704f7, 0xf9ba1651, 
	0x43103085, 0xfcdc1342, 0x48b2b335, 0xf69bf7c9, 0x4b418bbe, 0xf383a3e2, 0x45f704f7, 0xf9ba1651, 
	0x4fd288dc, 0xed6bf9d1, 0x4fd288dc, 0xed6bf9d1, 0x48b2b335, 0xf69bf7c9, 0x553805f2, 0xe4a2eff6, 
	0x539eba45, 0xe7821d59, 0x4b418bbe, 0xf383a3e2, 0x58c542c5, 0xdc71898d, 0x569cc31b, 0xe1d4a2c8, 
	0x4da1fab5, 0xf0730342, 0x5a6690ae, 0xd5052d97, 0x58c542c5, 0xdc71898d, 0x4fd288dc, 0xed6bf9d1, 
	0x5a12e720, 0xce86ff2a, 0x5a12e720, 0xd76619b6, 0x51d1dc80, 0xea70658a, 0x57cc15bc, 0xc91af976, 
	0x5a82799a, 0xd2bec333, 0x539eba45, 0xe7821d59, 0x539eba45, 0xc4df2862, 0x5a12e720, 0xce86ff2a, 
	0x553805f2, 0xe4a2eff6, 0x4da1fab5, 0xc1eb0209, 0x58c542c5, 0xcac933ae, 0x569cc31b, 0xe1d4a2c8, 
	0x45f704f7, 0xc04ee4b8, 0x569cc31b, 0xc78e9a1d, 0x57cc15bc, 0xdf18f0ce, 0x3cc85709, 0xc013bc39, 
	0x539eba45, 0xc4df2862, 0x58c542c5, 0xdc71898d, 0x3248d382, 0xc13ad060, 0x4fd288dc, 0xc2c17d52, 
	0x5987b08a, 0xd9e01006, 0x26b2a794, 0xc3bdbdf6, 0x4b418bbe, 0xc13ad060, 0x5a12e720, 0xd76619b6, 
	0x1a4608ab, 0xc78e9a1d, 0x45f704f7, 0xc04ee4b8, 0x5a6690ae, 0xd5052d97, 0x0d47d096, 0xcc983f70, 
	0x40000000, 0xc0000000, 0x5a82799a, 0xd2bec333, 0x00000000, 0xd2bec333, 0x396b3199, 0xc04ee4b8, 
	0x5a6690ae, 0xd09441bb, 0xf2b82f6a, 0xd9e01006, 0x3248d382, 0xc13ad060, 0x5a12e720, 0xce86ff2a, 
	0xe5b9f755, 0xe1d4a2c8, 0x2aaa7c7f, 0xc2c17d52, 0x5987b08a, 0xcc983f70, 0xd94d586c, 0xea70658a, 
	0x22a2f4f8, 0xc4df2862, 0x58c542c5, 0xcac933ae, 0xcdb72c7e, 0xf383a3e2, 0x1a4608ab, 0xc78e9a1d, 
	0x57cc15bc, 0xc91af976, 0xc337a8f7, 0xfcdc1342, 0x11a855df, 0xcac933ae, 0x569cc31b, 0xc78e9a1d, 
	0xba08fb09, 0x0645e9af, 0x08df1a8c, 0xce86ff2a, 0x553805f2, 0xc6250a18, 0xb25e054b, 0x0f8cfcbe, 
	0x00000000, 0xd2bec333, 0x539eba45, 0xc4df2862, 0xac6145bb, 0x187de2a7, 0xf720e574, 0xd76619b6, 
	0x51d1dc80, 0xc3bdbdf6, 0xa833ea44, 0x20e70f32, 0xee57aa21, 0xdc71898d, 0x4fd288dc, 0xc2c17d52, 
	0xa5ed18e0, 0x2899e64a, 0xe5b9f755, 0xe1d4a2c8, 0x4da1fab5, 0xc1eb0209, 0xa5996f52, 0x2f6bbe45, 
	0xdd5d0b08, 0xe7821d59, 0x4b418bbe, 0xc13ad060, 0xa73abd3b, 0x3536cc52, 0xd5558381, 0xed6bf9d1, 
	0x48b2b335, 0xc0b15502, 0xaac7fa0e, 0x39daf5e8, 0xcdb72c7e, 0xf383a3e2, 0x45f704f7, 0xc04ee4b8, 
	0xb02d7724, 0x3d3e82ae, 0xc694ce67, 0xf9ba1651, 0x43103085, 0xc013bc39, 0xb74d4ccb, 0x3f4eaafe, 
	
	0x40000000, 0x00000000, 0x40000000, 0x00000000, 0x40000000, 0x00000000, 0x418d2621, 0xfe6deaa1, 
	0x40c7d2bd, 0xff36f170, 0x424ff28f, 0xfda4f351, 0x43103085, 0xfcdc1342, 0x418d2621, 0xfe6deaa1, 
	0x4488e37f, 0xfb4ab7db, 0x4488e37f, 0xfb4ab7db, 0x424ff28f, 0xfda4f351, 0x46aa0d6d, 0xf8f21e8e, 
	0x45f704f7, 0xf9ba1651, 0x43103085, 0xfcdc1342, 0x48b2b335, 0xf69bf7c9, 0x475a5c77, 0xf82a6c6a, 
	0x43cdd89a, 0xfc135231, 0x4aa22036, 0xf4491311, 0x48b2b335, 0xf69bf7c9, 0x4488e37f, 0xfb4ab7db, 
	0x4c77a88e, 0xf1fa3ecb, 0x49ffd417, 0xf50ef5de, 0x454149fc, 0xfa824bfd, 0x4e32a956, 0xefb047f2, 
	0x4b418bbe, 0xf383a3e2, 0x45f704f7, 0xf9ba1651, 0x4fd288dc, 0xed6bf9d1, 0x4c77a88e, 0xf1fa3ecb, 
	0x46aa0d6d, 0xf8f21e8e, 0x5156b6d9, 0xeb2e1dbe, 0x4da1fab5, 0xf0730342, 0x475a5c77, 0xf82a6c6a, 
	0x52beac9f, 0xe8f77acf, 0x4ec05432, 0xeeee2d9d, 0x4807eb4b, 0xf7630799, 0x5409ed4b, 0xe6c8d59c, 
	0x4fd288dc, 0xed6bf9d1, 0x48b2b335, 0xf69bf7c9, 0x553805f2, 0xe4a2eff6, 0x50d86e6d, 0xebeca36c, 
	0x495aada2, 0xf5d544a7, 0x56488dc5, 0xe28688a4, 0x51d1dc80, 0xea70658a, 0x49ffd417, 0xf50ef5de, 
	0x573b2635, 0xe0745b24, 0x52beac9f, 0xe8f77acf, 0x4aa22036, 0xf4491311, 0x580f7b19, 0xde6d1f65, 
	0x539eba45, 0xe7821d59, 0x4b418bbe, 0xf383a3e2, 0x58c542c5, 0xdc71898d, 0x5471e2e6, 0xe61086bc, 
	0x4bde1089, 0xf2beafed, 0x595c3e2a, 0xda8249b4, 0x553805f2, 0xe4a2eff6, 0x4c77a88e, 0xf1fa3ecb, 
	0x59d438e5, 0xd8a00bae, 0x55f104dc, 0xe3399167, 0x4d0e4de2, 0xf136580d, 0x5a2d0957, 0xd6cb76c9, 
	0x569cc31b, 0xe1d4a2c8, 0x4da1fab5, 0xf0730342, 0x5a6690ae, 0xd5052d97, 0x573b2635, 0xe0745b24, 
	0x4e32a956, 0xefb047f2, 0x5a80baf6, 0xd34dcdb4, 0x57cc15bc, 0xdf18f0ce, 0x4ec05432, 0xeeee2d9d, 
	0x5a7b7f1a, 0xd1a5ef90, 0x584f7b58, 0xddc29958, 0x4f4af5d1, 0xee2cbbc1, 0x5a56deec, 0xd00e2639, 
	0x58c542c5, 0xdc71898d, 0x4fd288dc, 0xed6bf9d1, 0x5a12e720, 0xce86ff2a, 0x592d59da, 0xdb25f566, 
	0x50570819, 0xecabef3d, 0x59afaf4c, 0xcd110216, 0x5987b08a, 0xd9e01006, 0x50d86e6d, 0xebeca36c, 
	0x592d59da, 0xcbacb0bf, 0x59d438e5, 0xd8a00bae, 0x5156b6d9, 0xeb2e1dbe, 0x588c1404, 0xca5a86c4, 
	0x5a12e720, 0xd76619b6, 0x51d1dc80, 0xea70658a, 0x57cc15bc, 0xc91af976, 0x5a43b190, 0xd6326a88, 
	0x5249daa2, 0xe9b38223, 0x56eda1a0, 0xc7ee77b3, 0x5a6690ae, 0xd5052d97, 0x52beac9f, 0xe8f77acf, 
	0x55f104dc, 0xc6d569be, 0x5a7b7f1a, 0xd3de9156, 0x53304df6, 0xe83c56cf, 0x54d69714, 0xc5d03118, 
	0x5a82799a, 0xd2bec333, 0x539eba45, 0xe7821d59, 0x539eba45, 0xc4df2862, 0x5a7b7f1a, 0xd1a5ef90, 
	0x5409ed4b, 0xe6c8d59c, 0x5249daa2, 0xc402a33c, 0x5a6690ae, 0xd09441bb, 0x5471e2e6, 0xe61086bc, 
	0x50d86e6d, 0xc33aee27, 0x5a43b190, 0xcf89e3e8, 0x54d69714, 0xe55937d5, 0x4f4af5d1, 0xc2884e6e, 
	0x5a12e720, 0xce86ff2a, 0x553805f2, 0xe4a2eff6, 0x4da1fab5, 0xc1eb0209, 0x59d438e5, 0xcd8bbb6d, 
	0x55962bc0, 0xe3edb628, 0x4bde1089, 0xc1633f8a, 0x5987b08a, 0xcc983f70, 0x55f104dc, 0xe3399167, 
	0x49ffd417, 0xc0f1360b, 0x592d59da, 0xcbacb0bf, 0x56488dc5, 0xe28688a4, 0x4807eb4b, 0xc0950d1d, 
	0x58c542c5, 0xcac933ae, 0x569cc31b, 0xe1d4a2c8, 0x45f704f7, 0xc04ee4b8, 0x584f7b58, 0xc9edeb50, 
	0x56eda1a0, 0xe123e6ad, 0x43cdd89a, 0xc01ed535, 0x57cc15bc, 0xc91af976, 0x573b2635, 0xe0745b24, 
	0x418d2621, 0xc004ef3f, 0x573b2635, 0xc8507ea7, 0x57854ddd, 0xdfc606f1, 0x3f35b59d, 0xc0013bd3, 
	0x569cc31b, 0xc78e9a1d, 0x57cc15bc, 0xdf18f0ce, 0x3cc85709, 0xc013bc39, 0x55f104dc, 0xc6d569be, 
	0x580f7b19, 0xde6d1f65, 0x3a45e1f7, 0xc03c6a07, 0x553805f2, 0xc6250a18, 0x584f7b58, 0xddc29958, 
	0x37af354c, 0xc07b371e, 0x5471e2e6, 0xc57d965d, 0x588c1404, 0xdd196538, 0x350536f1, 0xc0d00db6, 
	0x539eba45, 0xc4df2862, 0x58c542c5, 0xdc71898d, 0x3248d382, 0xc13ad060, 0x52beac9f, 0xc449d892, 
	0x58fb0568, 0xdbcb0cce, 0x2f7afdfc, 0xc1bb5a11, 0x51d1dc80, 0xc3bdbdf6, 0x592d59da, 0xdb25f566, 
	0x2c9caf6c, 0xc2517e31, 0x50d86e6d, 0xc33aee27, 0x595c3e2a, 0xda8249b4, 0x29aee694, 0xc2fd08a9, 
	0x4fd288dc, 0xc2c17d52, 0x5987b08a, 0xd9e01006, 0x26b2a794, 0xc3bdbdf6, 0x4ec05432, 0xc2517e31, 
	0x59afaf4c, 0xd93f4e9e, 0x23a8fb93, 0xc4935b3c, 0x4da1fab5, 0xc1eb0209, 0x59d438e5, 0xd8a00bae, 
	0x2092f05f, 0xc57d965d, 0x4c77a88e, 0xc18e18a7, 0x59f54bee, 0xd8024d59, 0x1d719810, 0xc67c1e18, 
	0x4b418bbe, 0xc13ad060, 0x5a12e720, 0xd76619b6, 0x1a4608ab, 0xc78e9a1d, 0x49ffd417, 0xc0f1360b, 
	0x5a2d0957, 0xd6cb76c9, 0x17115bc0, 0xc8b4ab32, 0x48b2b335, 0xc0b15502, 0x5a43b190, 0xd6326a88, 
	0x13d4ae08, 0xc9edeb50, 0x475a5c77, 0xc07b371e, 0x5a56deec, 0xd59afadb, 0x10911f04, 0xcb39edca, 
	0x45f704f7, 0xc04ee4b8, 0x5a6690ae, 0xd5052d97, 0x0d47d096, 0xcc983f70, 0x4488e37f, 0xc02c64a6, 
	0x5a72c63b, 0xd4710883, 0x09f9e6a1, 0xce0866b8, 0x43103085, 0xc013bc39, 0x5a7b7f1a, 0xd3de9156, 
	0x06a886a0, 0xcf89e3e8, 0x418d2621, 0xc004ef3f, 0x5a80baf6, 0xd34dcdb4, 0x0354d741, 0xd11c3142, 
	0x40000000, 0xc0000000, 0x5a82799a, 0xd2bec333, 0x00000000, 0xd2bec333, 0x3e68fb62, 0xc004ef3f, 
	0x5a80baf6, 0xd2317756, 0xfcab28bf, 0xd4710883, 0x3cc85709, 0xc013bc39, 0x5a7b7f1a, 0xd1a5ef90, 
	0xf9577960, 0xd6326a88, 0x3b1e5335, 0xc02c64a6, 0x5a72c63b, 0xd11c3142, 0xf606195f, 0xd8024d59, 
	0x396b3199, 0xc04ee4b8, 0x5a6690ae, 0xd09441bb, 0xf2b82f6a, 0xd9e01006, 0x37af354c, 0xc07b371e, 
	0x5a56deec, 0xd00e2639, 0xef6ee0fc, 0xdbcb0cce, 0x35eaa2c7, 0xc0b15502, 0x5a43b190, 0xcf89e3e8, 
	0xec2b51f8, 0xddc29958, 0x341dbfd3, 0xc0f1360b, 0x5a2d0957, 0xcf077fe1, 0xe8eea440, 0xdfc606f1, 
	0x3248d382, 0xc13ad060, 0x5a12e720, 0xce86ff2a, 0xe5b9f755, 0xe1d4a2c8, 0x306c2624, 0xc18e18a7, 
	0x59f54bee, 0xce0866b8, 0xe28e67f0, 0xe3edb628, 0x2e88013a, 0xc1eb0209, 0x59d438e5, 0xcd8bbb6d, 
	0xdf6d0fa1, 0xe61086bc, 0x2c9caf6c, 0xc2517e31, 0x59afaf4c, 0xcd110216, 0xdc57046d, 0xe83c56cf, 
	0x2aaa7c7f, 0xc2c17d52, 0x5987b08a, 0xcc983f70, 0xd94d586c, 0xea70658a, 0x28b1b544, 0xc33aee27, 
	0x595c3e2a, 0xcc217822, 0xd651196c, 0xecabef3d, 0x26b2a794, 0xc3bdbdf6, 0x592d59da, 0xcbacb0bf, 
	0xd3635094, 0xeeee2d9d, 0x24ada23d, 0xc449d892, 0x58fb0568, 0xcb39edca, 0xd0850204, 0xf136580d, 
	0x22a2f4f8, 0xc4df2862, 0x58c542c5, 0xcac933ae, 0xcdb72c7e, 0xf383a3e2, 0x2092f05f, 0xc57d965d, 
	0x588c1404, 0xca5a86c4, 0xcafac90f, 0xf5d544a7, 0x1e7de5df, 0xc6250a18, 0x584f7b58, 0xc9edeb50, 
	0xc850cab4, 0xf82a6c6a, 0x1c6427a9, 0xc6d569be, 0x580f7b19, 0xc9836582, 0xc5ba1e09, 0xfa824bfd, 
	0x1a4608ab, 0xc78e9a1d, 0x57cc15bc, 0xc91af976, 0xc337a8f7, 0xfcdc1342, 0x1823dc7d, 0xc8507ea7, 
	0x57854ddd, 0xc8b4ab32, 0xc0ca4a63, 0xff36f170, 0x15fdf758, 0xc91af976, 0x573b2635, 0xc8507ea7, 
	0xbe72d9df, 0x0192155f, 0x13d4ae08, 0xc9edeb50, 0x56eda1a0, 0xc7ee77b3, 0xbc322766, 0x03ecadcf, 
	0x11a855df, 0xcac933ae, 0x569cc31b, 0xc78e9a1d, 0xba08fb09, 0x0645e9af, 0x0f7944a7, 0xcbacb0bf, 
	0x56488dc5, 0xc730e997, 0xb7f814b5, 0x089cf867, 0x0d47d096, 0xcc983f70, 0x55f104dc, 0xc6d569be, 
	0xb6002be9, 0x0af10a22, 0x0b145041, 0xcd8bbb6d, 0x55962bc0, 0xc67c1e18, 0xb421ef77, 0x0d415013, 
	0x08df1a8c, 0xce86ff2a, 0x553805f2, 0xc6250a18, 0xb25e054b, 0x0f8cfcbe, 0x06a886a0, 0xcf89e3e8, 
	0x54d69714, 0xc5d03118, 0xb0b50a2f, 0x11d3443f, 0x0470ebdc, 0xd09441bb, 0x5471e2e6, 0xc57d965d, 
	0xaf279193, 0x14135c94, 0x0238a1c6, 0xd1a5ef90, 0x5409ed4b, 0xc52d3d18, 0xadb6255e, 0x164c7ddd, 
	0x00000000, 0xd2bec333, 0x539eba45, 0xc4df2862, 0xac6145bb, 0x187de2a7, 0xfdc75e3a, 0xd3de9156, 
	0x53304df6, 0xc4935b3c, 0xab2968ec, 0x1aa6c82b, 0xfb8f1424, 0xd5052d97, 0x52beac9f, 0xc449d892, 
	0xaa0efb24, 0x1cc66e99, 0xf9577960, 0xd6326a88, 0x5249daa2, 0xc402a33c, 0xa9125e60, 0x1edc1953, 
	0xf720e574, 0xd76619b6, 0x51d1dc80, 0xc3bdbdf6, 0xa833ea44, 0x20e70f32, 0xf4ebafbf, 0xd8a00bae, 
	0x5156b6d9, 0xc37b2b6a, 0xa773ebfc, 0x22e69ac8, 0xf2b82f6a, 0xd9e01006, 0x50d86e6d, 0xc33aee27, 
	0xa6d2a626, 0x24da0a9a, 0xf086bb59, 0xdb25f566, 0x50570819, 0xc2fd08a9, 0xa65050b4, 0x26c0b162, 
	0xee57aa21, 0xdc71898d, 0x4fd288dc, 0xc2c17d52, 0xa5ed18e0, 0x2899e64a, 0xec2b51f8, 0xddc29958, 
	0x4f4af5d1, 0xc2884e6e, 0xa5a92114, 0x2a650525, 0xea0208a8, 0xdf18f0ce, 0x4ec05432, 0xc2517e31, 
	0xa58480e6, 0x2c216eaa, 0xe7dc2383, 0xe0745b24, 0x4e32a956, 0xc21d0eb8, 0xa57f450a, 0x2dce88aa, 
	0xe5b9f755, 0xe1d4a2c8, 0x4da1fab5, 0xc1eb0209, 0xa5996f52, 0x2f6bbe45, 0xe39bd857, 0xe3399167, 
	0x4d0e4de2, 0xc1bb5a11, 0xa5d2f6a9, 0x30f8801f, 0xe1821a21, 0xe4a2eff6, 0x4c77a88e, 0xc18e18a7, 
	0xa62bc71b, 0x32744493, 0xdf6d0fa1, 0xe61086bc, 0x4bde1089, 0xc1633f8a, 0xa6a3c1d6, 0x33de87de, 
	0xdd5d0b08, 0xe7821d59, 0x4b418bbe, 0xc13ad060, 0xa73abd3b, 0x3536cc52, 0xdb525dc3, 0xe8f77acf, 
	0x4aa22036, 0xc114ccb9, 0xa7f084e7, 0x367c9a7e, 0xd94d586c, 0xea70658a, 0x49ffd417, 0xc0f1360b, 
	0xa8c4d9cb, 0x37af8159, 0xd74e4abc, 0xebeca36c, 0x495aada2, 0xc0d00db6, 0xa9b7723b, 0x38cf1669, 
	0xd5558381, 0xed6bf9d1, 0x48b2b335, 0xc0b15502, 0xaac7fa0e, 0x39daf5e8, 0xd3635094, 0xeeee2d9d, 
	0x4807eb4b, 0xc0950d1d, 0xabf612b5, 0x3ad2c2e8, 0xd177fec6, 0xf0730342, 0x475a5c77, 0xc07b371e, 
	0xad415361, 0x3bb6276e, 0xcf93d9dc, 0xf1fa3ecb, 0x46aa0d6d, 0xc063d405, 0xaea94927, 0x3c84d496, 
	0xcdb72c7e, 0xf383a3e2, 0x45f704f7, 0xc04ee4b8, 0xb02d7724, 0x3d3e82ae, 0xcbe2402d, 0xf50ef5de, 
	0x454149fc, 0xc03c6a07, 0xb1cd56aa, 0x3de2f148, 0xca155d39, 0xf69bf7c9, 0x4488e37f, 0xc02c64a6, 
	0xb3885772, 0x3e71e759, 0xc850cab4, 0xf82a6c6a, 0x43cdd89a, 0xc01ed535, 0xb55ddfca, 0x3eeb3347, 
	0xc694ce67, 0xf9ba1651, 0x43103085, 0xc013bc39, 0xb74d4ccb, 0x3f4eaafe, 0xc4e1accb, 0xfb4ab7db, 
	0x424ff28f, 0xc00b1a20, 0xb955f293, 0x3f9c2bfb, 0xc337a8f7, 0xfcdc1342, 0x418d2621, 0xc004ef3f, 
	0xbb771c81, 0x3fd39b5a, 0xc197049e, 0xfe6deaa1, 0x40c7d2bd, 0xc0013bd3, 0xbdb00d71, 0x3ff4e5e0, 
};
*/
