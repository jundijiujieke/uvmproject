module imdct_rom576x64(
clk,
en,
addr,

dout
);

input clk;
input en;
input [9:0] addr;

output reg [63:0] dout;

reg [63:0] mem[0:575]={ 

64'hbf9bc731_ff9b783c, 
64'hbed5332c_c002c697,
64'hbe112251_fe096c8d,
64'hbd4f9c30_c00f1c4a, 
64'hbc90a83f_fc77ae5e, 
64'hbbd44dd9_c0254e27, 
64'hbb1a9443_fae67ba2, 
64'hba6382a6_c04558c0, 
64'hb9af200f_f9561237, 
64'hb8fd7373_c06f3726, 
64'hb84e83ac_f7c6afdc, 
64'hb7a25779_c0a2e2e3, 
64'hb6f8f57c_f6389228, 
64'hb652643e_c0e05401, 
64'hb5aeaa2a_f4abf67e, 
64'hb50dcd90_c1278104, 
64'hb46fd4a4_f3211a07, 
64'hb3d4c57c_c1785ef4, 
64'hb33ca614_f19839a6, 
64'hb2a77c49_c1d2e158, 
64'hb2154dda_f01191f3, 
64'hb186206b_c236fa3b, 
64'hb0f9f981_ee8d5f29, 
64'hb070de82_c2a49a2e, 
64'hafead4b9_ed0bdd25, 
64'haf67e14f_c31bb049, 
64'haee80952_eb8d475b, 
64'hae6b51ae_c39c2a2f, 
64'hadf1bf34_ea11d8c8, 
64'had7b5692_c425f410, 
64'had081c5a_e899cbf1, 
64'hac9814fd_c4b8f8ad, 
64'hac2b44cc_e7255ad1, 
64'habc1aff9_c555215a, 
64'hab5b5a96_e5b4bed8, 
64'haaf84896_c5fa5603, 
64'haa987dca_e44830dd, 
64'haa3bfde3_c6a87d2d, 
64'ha9e2cc73_e2dfe917, 
64'ha98cece9_c75f7bfe, 
64'ha93a6296_e17c1f15, 
64'ha8eb30a7_c81f363d, 
64'ha89f5a2b_e01d09b4, 
64'ha856e20e_c8e78e5b, 
64'ha811cb1b_dec2df18, 
64'ha7d017fc_c9b86572, 
64'ha791cb39_dd6dd4a2, 
64'ha756e73a_ca919b4e, 
64'ha71f6e43_dc1e1ee9, 
64'ha6eb6279_cb730e70, 
64'ha6bac5dc_dad3f1b1, 
64'ha68d9a4c_cc5c9c14, 
64'ha663e188_d98f7fe6, 
64'ha63d9d2b_cd4e2037, 
64'ha61aceaf_d850fb8e, 
64'ha5fb776b_ce47759a, 
64'ha5df9894_d71895c9, 
64'ha5c7333e_cf4875ca, 
64'ha5b2485a_d5e67ec1, 
64'ha5a0d8b5_d050f926, 
64'ha592e4fd_d4bae5ab, 
64'ha5886dba_d160d6e5, 
64'ha5817354_d395f8ba, 
64'ha57df60f_d277e518, 
/* 1024 - format = Q30 * 2^-10 */
64'hbff3703e_fff36f02, 
64'hbfda5824_c0000b1a, 
64'hbfc149ed_ffc12b16, 
64'hbfa845a0_c0003c74, 
64'hbf8f4b3e_ff8ee750, 
64'hbf765acc_c0009547, 
64'hbf5d744e_ff5ca3d0, 
64'hbf4497c8_c0011594, 
64'hbf2bc53d_ff2a60b4, 
64'hbf12fcb2_c001bd5c, 
64'hbefa3e2a_fef81e1d, 
64'hbee189a8_c0028c9c, 
64'hbec8df32_fec5dc28, 
64'hbeb03eca_c0038356, 
64'hbe97a875_fe939af5, 
64'hbe7f1c36_c004a188, 
64'hbe669a10_fe615aa3, 
64'hbe4e2209_c005e731, 
64'hbe35b423_fe2f1b50, 
64'hbe1d5062_c0075452, 
64'hbe04f6cb_fdfcdd1d, 
64'hbdeca760_c008e8e8, 
64'hbdd46225_fdcaa027, 
64'hbdbc2720_c00aa4f3, 
64'hbda3f652_fd98648d, 
64'hbd8bcfbf_c00c8872, 
64'hbd73b36d_fd662a70, 
64'hbd5ba15d_c00e9364, 
64'hbd439995_fd33f1ed, 
64'hbd2b9c17_c010c5c7, 
64'hbd13a8e7_fd01bb24, 
64'hbcfbc00a_c0131f9b, 
64'hbce3e182_fccf8634, 
64'hbccc0d53_c015a0dd, 
64'hbcb44382_fc9d533b, 
64'hbc9c8411_c018498c, 
64'hbc84cf05_fc6b2259, 
64'hbc6d2461_c01b19a7, 
64'hbc558428_fc38f3ac, 
64'hbc3dee5f_c01e112b, 
64'hbc266309_fc06c754, 
64'hbc0ee22a_c0213018, 
64'hbbf76bc4_fbd49d70, 
64'hbbdfffdd_c024766a, 
64'hbbc89e77_fba2761e, 
64'hbbb14796_c027e421, 
64'hbb99fb3e_fb70517d, 
64'hbb82b972_c02b7939, 
64'hbb6b8235_fb3e2fac, 
64'hbb54558d_c02f35b1, 
64'hbb3d337b_fb0c10cb, 
64'hbb261c04_c0331986, 
64'hbb0f0f2b_fad9f4f8, 
64'hbaf80cf4_c03724b6, 
64'hbae11561_faa7dc52, 
64'hbaca2878_c03b573f, 
64'hbab3463b_fa75c6f8, 
64'hba9c6eae_c03fb11d, 
64'hba85a1d4_fa43b508, 
64'hba6edfb1_c044324f, 
64'hba582849_fa11a6a3, 
64'hba417b9e_c048dad1, 
64'hba2ad9b5_f9df9be6, 
64'hba144291_c04daaa1, 
64'hb9fdb635_f9ad94f0, 
64'hb9e734a4_c052a1bb, 
64'hb9d0bde4_f97b91e1, 
64'hb9ba51f6_c057c01d, 
64'hb9a3f0de_f94992d7, 
64'hb98d9aa0_c05d05c3, 
64'hb9774f3f_f91797f0, 
64'hb9610ebe_c06272aa, 
64'hb94ad922_f8e5a14d, 
64'hb934ae6d_c06806ce, 
64'hb91e8ea3_f8b3af0c, 
64'hb90879c7_c06dc22e, 
64'hb8f26fdc_f881c14b, 
64'hb8dc70e7_c073a4c3, 
64'hb8c67cea_f84fd829, 
64'hb8b093ea_c079ae8c, 
64'hb89ab5e8_f81df3c5, 
64'hb884e2e9_c07fdf85, 
64'hb86f1af0_f7ec143e, 
64'hb8595e00_c08637a9, 
64'hb843ac1d_f7ba39b3, 
64'hb82e0549_c08cb6f5, 
64'hb818698a_f7886442, 
64'hb802d8e0_c0935d64, 
64'hb7ed5351_f756940a, 
64'hb7d7d8df_c09a2af3, 
64'hb7c2698e_f724c92a, 
64'hb7ad0561_c0a11f9d, 
64'hb797ac5b_f6f303c0, 
64'hb7825e80_c0a83b5e, 
64'hb76d1bd2_f6c143ec, 
64'hb757e455_c0af7e33, 
64'hb742b80d_f68f89cb, 
64'hb72d96fd_c0b6e815, 
64'hb7188127_f65dd57d, 
64'hb7037690_c0be7901, 
64'hb6ee773a_f62c2721, 
64'hb6d98328_c0c630f2, 
64'hb6c49a5e_f5fa7ed4, 
64'hb6afbce0_c0ce0fe3, 
64'hb69aeab0_f5c8dcb6, 
64'hb68623d1_c0d615cf, 
64'hb6716847_f59740e5, 
64'hb65cb815_c0de42b2, 
64'hb648133e_f565ab80, 
64'hb63379c5_c0e69686, 
64'hb61eebae_f5341ca5, 
64'hb60a68fb_c0ef1147, 
64'hb5f5f1b1_f5029473, 
64'hb5e185d1_c0f7b2ee, 
64'hb5cd255f_f4d11308, 
64'hb5b8d05f_c1007b77, 
64'hb5a486d2_f49f9884, 
64'hb59048be_c1096add, 
64'hb57c1624_f46e2504, 
64'hb567ef08_c1128119, 
64'hb553d36c_f43cb8a7, 
64'hb53fc355_c11bbe26, 
64'hb52bbec4_f40b538b, 
64'hb517c5be_c12521ff, 
64'hb503d845_f3d9f5cf, 
64'hb4eff65c_c12eac9d, 
64'hb4dc2007_f3a89f92, 
64'hb4c85548_c1385dfb, 
64'hb4b49622_f37750f2, 
64'hb4a0e299_c1423613, 
64'hb48d3ab0_f3460a0d, 
64'hb4799e69_c14c34df, 
64'hb4660dc8_f314cb02, 
64'hb45288cf_c1565a58, 
64'hb43f0f82_f2e393ef, 
64'hb42ba1e4_c160a678, 
64'hb4183ff7_f2b264f2, 
64'hb404e9bf_c16b193a, 
64'hb3f19f3e_f2813e2a, 
64'hb3de6078_c175b296, 
64'hb3cb2d70_f2501fb5, 
64'hb3b80628_c1807285, 
64'hb3a4eaa4_f21f09b1, 
64'hb391dae6_c18b5903, 
64'hb37ed6f1_f1edfc3d, 
64'hb36bdec9_c1966606, 
64'hb358f26f_f1bcf777, 
64'hb34611e8_c1a1998a, 
64'hb3333d36_f18bfb7d, 
64'hb320745c_c1acf386, 
64'hb30db75d_f15b086d, 
64'hb2fb063b_c1b873f5, 
64'hb2e860fa_f12a1e66, 
64'hb2d5c79d_c1c41ace, 
64'hb2c33a26_f0f93d86, 
64'hb2b0b898_c1cfe80a, 
64'hb29e42f6_f0c865ea, 
64'hb28bd943_c1dbdba3, 
64'hb2797b82_f09797b2, 
64'hb26729b5_c1e7f591, 
64'hb254e3e0_f066d2fa, 
64'hb242aa05_c1f435cc, 
64'hb2307c27_f03617e2, 
64'hb21e5a49_c2009c4e, 
64'hb20c446d_f0056687, 
64'hb1fa3a97_c20d290d, 
64'hb1e83cc9_efd4bf08, 
64'hb1d64b06_c219dc03, 
64'hb1c46551_efa42181, 
64'hb1b28bad_c226b528, 
64'hb1a0be1b_ef738e12, 
64'hb18efca0_c233b473, 
64'hb17d473d_ef4304d8, 
64'hb16b9df6_c240d9de, 
64'hb15a00cd_ef1285f2, 
64'hb1486fc5_c24e255e, 
64'hb136eae1_eee2117c, 
64'hb1257223_c25b96ee, 
64'hb114058e_eeb1a796, 
64'hb102a524_c2692e83, 
64'hb0f150e9_ee81485c, 
64'hb0e008e0_c276ec16, 
64'hb0cecd09_ee50f3ed, 
64'hb0bd9d6a_c284cf9f, 
64'hb0ac7a03_ee20aa67, 
64'hb09b62d8_c292d914, 
64'hb08a57eb_edf06be6, 
64'hb079593f_c2a1086d, 
64'hb06866d7_edc0388a, 
64'hb05780b5_c2af5da2, 
64'hb046a6db_ed901070, 
64'hb035d94e_c2bdd8a9, 
64'hb025180e_ed5ff3b5, 
64'hb014631e_c2cc7979, 
64'hb003ba82_ed2fe277, 
64'haff31e3b_c2db400a, 
64'hafe28e4d_ecffdcd4, 
64'hafd20ab9_c2ea2c53, 
64'hafc19383_eccfe2ea, 
64'hafb128ad_c2f93e4a, 
64'hafa0ca39_ec9ff4d6, 
64'haf90782a_c30875e5, 
64'haf803283_ec7012b5, 
64'haf6ff945_c317d31c, 
64'haf5fcc74_ec403ca5, 
64'haf4fac12_c32755e5, 
64'haf3f9822_ec1072c4, 
64'haf2f90a5_c336fe37, 
64'haf1f959f_ebe0b52f, 
64'haf0fa712_c346cc07, 
64'haeffc500_ebb10404, 
64'haeefef6c_c356bf4d, 
64'haee02658_eb815f60, 
64'haed069c7_c366d7fd, 
64'haec0b9bb_eb51c760, 
64'haeb11636_c377160f, 
64'haea17f3b_eb223c22, 
64'hae91f4cd_c3877978, 
64'hae8276ed_eaf2bdc3, 
64'hae73059f_c398022f, 
64'hae63a0e3_eac34c60, 
64'hae5448be_c3a8b028, 
64'hae44fd31_ea93e817, 
64'hae35be3f_c3b9835a, 
64'hae268be9_ea649105, 
64'hae176633_c3ca7bba, 
64'hae084d1f_ea354746, 
64'hadf940ae_c3db993e, 
64'hadea40e4_ea060af9, 
64'haddb4dc2_c3ecdbdc, 
64'hadcc674b_e9d6dc3b, 
64'hadbd8d82_c3fe4388, 
64'hadaec067_e9a7bb28, 
64'had9fffff_c40fd037, 
64'had914c4b_e978a7dd, 
64'had82a54c_c42181e0, 
64'had740b07_e949a278, 
64'had657d7c_c4335877, 
64'had56fcaf_e91aab16, 
64'had4888a0_c44553f2, 
64'had3a2153_e8ebc1d3, 
64'had2bc6ca_c4577444, 
64'had1d7907_e8bce6cd, 
64'had0f380c_c469b963, 
64'had0103db_e88e1a20, 
64'hacf2dc77_c47c2344, 
64'hace4c1e2_e85f5be9, 
64'hacd6b41e_c48eb1db, 
64'hacc8b32c_e830ac45, 
64'hacbabf10_c4a1651c, 
64'hacacd7cb_e8020b52, 
64'hac9efd60_c4b43cfd, 
64'hac912fd1_e7d3792b, 
64'hac836f1f_c4c73972, 
64'hac75bb4d_e7a4f5ed, 
64'hac68145d_c4da5a6f, 
64'hac5a7a52_e77681b6, 
64'hac4ced2c_c4ed9fe7, 
64'hac3f6cef_e7481ca1, 
64'hac31f99d_c50109d0, 
64'hac249336_e719c6cb, 
64'hac1739bf_c514981d, 
64'hac09ed38_e6eb8052, 
64'habfcada3_c5284ac3, 
64'habef7b04_e6bd4951, 
64'habe2555b_c53c21b4, 
64'habd53caa_e68f21e5, 
64'habc830f5_c5501ce5, 
64'habbb323c_e6610a2a, 
64'habae4082_c5643c4a, 
64'haba15bc9_e633023e, 
64'hab948413_c5787fd6, 
64'hab87b962_e6050a3b, 
64'hab7afbb7_c58ce77c, 
64'hab6e4b15_e5d72240, 
64'hab61a77d_c5a17330, 
64'hab5510f3_e5a94a67, 
64'hab488776_c5b622e6, 
64'hab3c0b0b_e57b82cd, 
64'hab2f9bb1_c5caf690, 
64'hab23396c_e54dcb8f, 
64'hab16e43d_c5dfee22, 
64'hab0a9c27_e52024c9, 
64'haafe612a_c5f5098f, 
64'haaf23349_e4f28e96, 
64'haae61286_c60a48c9, 
64'haad9fee3_e4c50914, 
64'haacdf861_c61fabc4, 
64'haac1ff03_e497945d, 
64'haab612ca_c6353273, 
64'haaaa33b8_e46a308f, 
64'haa9e61cf_c64adcc7, 
64'haa929d10_e43cddc4, 
64'haa86e57e_c660aab5, 
64'haa7b3b1b_e40f9c1a, 
64'haa6f9de7_c6769c2e, 
64'haa640de6_e3e26bac, 
64'haa588b18_c68cb124, 
64'haa4d157f_e3b54c95, 
64'haa41ad1e_c6a2e98b, 
64'haa3651f6_e3883ef2, 
64'haa2b0409_c6b94554, 
64'haa1fc358_e35b42df, 
64'haa148fe6_c6cfc472, 
64'haa0969b3_e32e5876, 
64'ha9fe50c2_c6e666d7, 
64'ha9f34515_e3017fd5, 
64'ha9e846ad_c6fd2c75, 
64'ha9dd558b_e2d4b916, 
64'ha9d271b2_c714153e, 
64'ha9c79b23_e2a80456, 
64'ha9bcd1e0_c72b2123, 
64'ha9b215ea_e27b61af, 
64'ha9a76744_c7425016, 
64'ha99cc5ee_e24ed13d, 
64'ha99231eb_c759a20a, 
64'ha987ab3c_e222531c, 
64'ha97d31e3_c77116f0, 
64'ha972c5e1_e1f5e768, 
64'ha9686738_c788aeb9, 
64'ha95e15e9_e1c98e3b, 
64'ha953d1f7_c7a06957, 
64'ha9499b62_e19d47b1, 
64'ha93f722c_c7b846ba, 
64'ha9355658_e17113e5, 
64'ha92b47e5_c7d046d6, 
64'ha92146d7_e144f2f3, 
64'ha917532e_c7e8699a, 
64'ha90d6cec_e118e4f6, 
64'ha9039413_c800aef7, 
64'ha8f9c8a4_e0ecea09, 
64'ha8f00aa0_c81916df, 
64'ha8e65a0a_e0c10247, 
64'ha8dcb6e2_c831a143, 
64'ha8d3212a_e0952dcb, 
64'ha8c998e3_c84a4e14, 
64'ha8c01e10_e0696cb0, 
64'ha8b6b0b1_c8631d42, 
64'ha8ad50c8_e03dbf11, 
64'ha8a3fe57_c87c0ebd, 
64'ha89ab95e_e012250a, 
64'ha89181df_c8952278, 
64'ha88857dc_dfe69eb4, 
64'ha87f3b57_c8ae5862, 
64'ha8762c4f_dfbb2c2c, 
64'ha86d2ac8_c8c7b06b, 
64'ha86436c2_df8fcd8b, 
64'ha85b503e_c8e12a84, 
64'ha852773f_df6482ed, 
64'ha849abc4_c8fac69e, 
64'ha840edd1_df394c6b, 
64'ha8383d66_c91484a8, 
64'ha82f9a84_df0e2a22, 
64'ha827052d_c92e6492, 
64'ha81e7d62_dee31c2b, 
64'ha8160324_c948664d, 
64'ha80d9675_deb822a1, 
64'ha8053756_c96289c9, 
64'ha7fce5c9_de8d3d9e, 
64'ha7f4a1ce_c97ccef5, 
64'ha7ec6b66_de626d3e, 
64'ha7e44294_c99735c2, 
64'ha7dc2759_de37b199, 
64'ha7d419b4_c9b1be1e, 
64'ha7cc19a9_de0d0acc, 
64'ha7c42738_c9cc67fa, 
64'ha7bc4262_dde278ef, 
64'ha7b46b29_c9e73346, 
64'ha7aca18e_ddb7fc1e, 
64'ha7a4e591_ca021fef, 
64'ha79d3735_dd8d9472, 
64'ha795967a_ca1d2de7, 
64'ha78e0361_dd634206, 
64'ha7867dec_ca385d1d, 
64'ha77f061c_dd3904f4, 
64'ha7779bf2_ca53ad7e, 
64'ha7703f70_dd0edd55, 
64'ha768f095_ca6f1efc, 
64'ha761af64_dce4cb44, 
64'ha75a7bdd_ca8ab184, 
64'ha7535602_dcbacedb, 
64'ha74c3dd4_caa66506, 
64'ha7453353_dc90e834, 
64'ha73e3681_cac23971, 
64'ha7374760_dc671768, 
64'ha73065ef_cade2eb3, 
64'ha7299231_dc3d5c91, 
64'ha722cc25_cafa44bc, 
64'ha71c13ce_dc13b7c9, 
64'ha715692c_cb167b79, 
64'ha70ecc41_dbea292b, 
64'ha7083d0d_cb32d2da, 
64'ha701bb91_dbc0b0ce, 
64'ha6fb47ce_cb4f4acd, 
64'ha6f4e1c6_db974ece, 
64'ha6ee8979_cb6be341, 
64'ha6e83ee8_db6e0342, 
64'ha6e20214_cb889c23, 
64'ha6dbd2ff_db44ce46, 
64'ha6d5b1a9_cba57563, 
64'ha6cf9e13_db1baff2, 
64'ha6c9983e_cbc26eee, 
64'ha6c3a02b_daf2a860, 
64'ha6bdb5da_cbdf88b3, 
64'ha6b7d94e_dac9b7a9, 
64'ha6b20a86_cbfcc29f, 
64'ha6ac4984_daa0dde7, 
64'ha6a69649_cc1a1ca0, 
64'ha6a0f0d5_da781b31, 
64'ha69b5929_cc3796a5, 
64'ha695cf46_da4f6fa3, 
64'ha690532d_cc55309b, 
64'ha68ae4df_da26db54, 
64'ha685845c_cc72ea70, 
64'ha68031a6_d9fe5e5e, 
64'ha67aecbd_cc90c412, 
64'ha675b5a3_d9d5f8d9, 
64'ha6708c57_ccaebd6e, 
64'ha66b70db_d9adaadf, 
64'ha6666330_ccccd671, 
64'ha6616355_d9857489, 
64'ha65c714d_cceb0f0a, 
64'ha6578d18_d95d55ef, 
64'ha652b6b6_cd096725, 
64'ha64dee28_d9354f2a, 
64'ha6493370_cd27deb0, 
64'ha644868d_d90d6053, 
64'ha63fe781_cd467599, 
64'ha63b564c_d8e58982, 
64'ha636d2ee_cd652bcb, 
64'ha6325d6a_d8bdcad0, 
64'ha62df5bf_cd840134, 
64'ha6299bed_d8962456, 
64'ha6254ff7_cda2f5c2, 
64'ha62111db_d86e962b, 
64'ha61ce19c_cdc20960, 
64'ha618bf39_d8472069, 
64'ha614aab3_cde13bfd, 
64'ha610a40c_d81fc328, 
64'ha60cab43_ce008d84, 
64'ha608c058_d7f87e7f, 
64'ha604e34e_ce1ffde2, 
64'ha6011424_d7d15288, 
64'ha5fd52db_ce3f8d05, 
64'ha5f99f73_d7aa3f5a, 
64'ha5f5f9ed_ce5f3ad8, 
64'ha5f2624a_d783450d, 
64'ha5eed88a_ce7f0748, 
64'ha5eb5cae_d75c63ba, 
64'ha5e7eeb6_ce9ef241, 
64'ha5e48ea3_d7359b78, 
64'ha5e13c75_cebefbb0, 
64'ha5ddf82d_d70eec60, 
64'ha5dac1cb_cedf2380, 
64'ha5d79950_d6e85689, 
64'ha5d47ebc_ceff699f, 
64'ha5d17210_d6c1da0b, 
64'ha5ce734d_cf1fcdf8, 
64'ha5cb8272_d69b76fe, 
64'ha5c89f80_cf405077, 
64'ha5c5ca77_d6752d79, 
64'ha5c30359_cf60f108, 
64'ha5c04a25_d64efd94, 
64'ha5bd9edc_cf81af97, 
64'ha5bb017f_d628e767, 
64'ha5b8720d_cfa28c10, 
64'ha5b5f087_d602eb0a, 
64'ha5b37cee_cfc3865e, 
64'ha5b11741_d5dd0892, 
64'ha5aebf82_cfe49e6d, 
64'ha5ac75b0_d5b74019, 
64'ha5aa39cd_d005d42a, 
64'ha5a80bd7_d59191b5, 
64'ha5a5ebd0_d027277e, 
64'ha5a3d9b8_d56bfd7d, 
64'ha5a1d590_d0489856, 
64'ha59fdf57_d5468389, 
64'ha59df70e_d06a269d, 
64'ha59c1cb5_d52123f0, 
64'ha59a504c_d08bd23f, 
64'ha59891d4_d4fbdec9, 
64'ha596e14e_d0ad9b26, 
64'ha5953eb8_d4d6b42b, 
64'ha593aa14_d0cf813e, 
64'ha5922362_d4b1a42c, 
64'ha590aaa2_d0f18472, 
64'ha58f3fd4_d48caee4, 
64'ha58de2f8_d113a4ad, 
64'ha58c940f_d467d469, 
64'ha58b5319_d135e1d9, 
64'ha58a2016_d44314d3, 
64'ha588fb06_d1583be2, 
64'ha587e3ea_d41e7037, 
64'ha586dac1_d17ab2b3, 
64'ha585df8c_d3f9e6ad, 
64'ha584f24b_d19d4636, 
64'ha58412fe_d3d5784a, 
64'ha58341a5_d1bff656, 
64'ha5827e40_d3b12526, 
64'ha581c8d0_d1e2c2fd, 
64'ha5812154_d38ced57, 
64'ha58087cd_d205ac17, 
64'ha57ffc3b_d368d0f3, 
64'ha57f7e9d_d228b18d, 
64'ha57f0ef5_d344d011, 
64'ha57ead41_d24bd34a, 
64'ha57e5982_d320eac6, 
64'ha57e13b8_d26f1138, 
64'ha57ddbe4_d2fd2129, 
64'ha57db204_d2926b41, 
64'ha57d961a_d2d97350, 
64'ha57d8825_d2b5e151 
};


always @(posedge clk) 
  if (en)
    dout <= mem[addr];

endmodule
